module CUT (GND,VDD,CK,SE,SI,SO,g100,g101,g102,g103,g10377,g10379,g104,g10455,g10457,g10459,g10461,g10463,g10465,g10628,g10801,g109,g11163,g11206,g11489,g1170,g1173,g1176,g1179,g1182,g1185,g1188,g1191,g1194,g1197,g1200,g1203,g1696,g1700,g1712,g18,g1957,g1960,g1961,g23,g2355,g2601,g2602,g2603,g2604,g2605,g2606,g2607,g2608,g2609,g2610,g2611,g2612,g2648,g27,g28,g29,g2986,g30,g3007,g3069,g31,g3327,g41,g4171,g4172,g4173,g4174,g4175,g4176,g4177,g4178,g4179,g4180,g4181,g4191,g4192,g4193,g4194,g4195,g4196,g4197,g4198,g4199,g42,g4200,g4201,g4202,g4203,g4204,g4205,g4206,g4207,g4208,g4209,g4210,g4211,g4212,g4213,g4214,g4215,g4216,g43,g44,g45,g46,g47,g48,g4887,g4888,g5101,g5105,g5658,g5659,g5816,g6253,g6254,g6255,g6256,g6257,g6258,g6259,g6260,g6261,g6262,g6263,g6264,g6265,g6266,g6267,g6268,g6269,g6270,g6271,g6272,g6273,g6274,g6275,g6276,g6277,g6278,g6279,g6280,g6281,g6282,g6283,g6284,g6285,g6842,g6920,g6926,g6932,g6942,g6949,g6955,g741,g742,g743,g744,g750,g7744,g8061,g8062,g82,g8271,g83,g8313,g8316,g8318,g8323,g8328,g8331,g8335,g8340,g8347,g8349,g8352,g84,g85,g8561,g8562,g8563,g8564,g8565,g8566,g86,g87,g872,g873,g877,g88,g881,g886,g889,g89,g892,g895,g8976,g8977,g8978,g8979,g898,g8980,g8981,g8982,g8983,g8984,g8985,g8986,g90,g901,g904,g907,g91,g910,g913,g916,g919,g92,g922,g925,g93,g94,g9451,g95,g96,g99,g9961);
input GND,VDD,CK,SE,SI,g18,g27,g109,g741,g742,g743,g744,g872,g873,g877,g881,g1712,g1960,g1961,g1696,g750,g85,g42,g1700,g102,g104,g101,g29,g28,g103,g83,g23,g87,g922,g892,g84,g919,g1182,g925,g48,g895,g889,g1185,g41,g43,g99,g1173,g1203,g1188,g1197,g46,g31,g45,g92,g89,g898,g91,g93,g913,g82,g88,g1194,g47,g96,g910,g95,g904,g1176,g901,g44,g916,g100,g886,g30,g86,g1170,g1200,g1191,g907,g90,g94,g1179;
output SO,g2355,g2601,g2602,g2603,g2604,g2605,g2606,g2607,g2608,g2609,g2610,g2611,g2612,g2648,g2986,g3007,g3069,g4172,g4173,g4174,g4175,g4176,g4177,g4178,g4179,g4180,g4181,g4887,g4888,g5101,g5105,g5658,g5659,g5816,g6920,g6926,g6932,g6942,g6949,g6955,g7744,g8061,g8062,g8271,g8313,g8316,g8318,g8323,g8328,g8331,g8335,g8340,g8347,g8349,g8352,g8561,g8562,g8563,g8564,g8565,g8566,g8976,g8977,g8978,g8979,g8980,g8981,g8982,g8983,g8984,g8985,g8986,g9451,g9961,g10377,g10379,g10455,g10457,g10459,g10461,g10463,g10465,g10628,g10801,g11163,g11206,g11489,g6842,g4171,g6267,g6257,g1957,g6282,g6284,g6281,g6253,g6285,g6283,g6265,g3327,g6269,g4204,g4193,g6266,g4203,g4212,g4196,g6263,g4194,g4192,g4213,g6256,g6258,g6279,g4209,g4208,g4214,g4206,g6261,g6255,g6260,g6274,g6271,g4195,g6273,g6275,g4201,g6264,g6270,g4216,g6262,g6278,g4200,g6277,g4198,g4210,g4197,g6259,g4202,g6280,g4191,g6254,g6268,g4205,g4207,g4215,g4199,g6272,g6276,g4211;
wire SE_B,CK1,CK2,g1289,g5660,g1882,g9349,g312,g5644,g452,g11257,g123,g8272,g207,g7315,g713,g9345,g1153,g6304,g1209,g10873,g1744,g5663,g1558,g7349,g695,g9343,g461,g11467,g940,g8572,g976,g11471,g709,g8432,g1092,g6810,g1574,g7354,g1864,g7816,g369,g11439,g1580,g7356,g1736,g6846,g39,g10774,g1651,g11182,g1424,g7330,g1737,g1672,g11037,g1077,g6805,g1231,g8279,g4,g8079,g774,g7785,g1104,g6815,g1304,g7290,g243,g7325,g1499,g8447,g1044,g7789,g1444,g8987,g757,g11179,g786,g8436,g1543,g7344,g552,g11045,g315,g5645,g1534,g7341,g622,g9338,g1927,g9354,g1660,g11033,g278,g7765,g1436,g8989,g718,g8433,g76,g7775,g554,g11047,g496,g11333,g981,g11472,g878,g4896,g590,g5653,g829,g4182,g1095,g6811,g704,g9344,g1265,g7302,g1786,g7814,g682,g8429,g1296,g7292,g587,g6295,g52,g7777,g646,g8065,g327,g5649,g1389,g6836,g1371,g7311,g1956,g1955,g1675,g11038,g354,g11508,g113,g7285,g639,g8063,g1684,g11041,g1639,g8448,g1791,g8080,g248,g7323,g1707,g4907,g1759,g5668,g351,g11507,g1604,g7364,g1098,g6812,g932,g8570,g126,g5642,g1896,g8282,g736,g8435,g1019,g7807,g1362,g7305,g745,g2639,g1419,g7332,g58,g7779,g32,g11397,g876,g1086,g6808,g1486,g8444,g1730,g10881,g1504,g7328,g1470,g8440,g822,g8437,g583,g6291,g1678,g11039,g174,g8423,g1766,g7810,g1801,g8450,g186,g7317,g959,g11403,g1169,g6314,g1007,g7806,g1407,g8993,g1059,g7794,g1868,g7817,g758,g6797,g1718,g6337,g396,g11265,g1015,g7808,g38,g10872,g632,g5655,g1415,g7335,g1227,g8278,g1721,g10878,g882,g883,g16,g4906,g284,g7767,g426,g11256,g219,g7310,g1216,g1360,g806,g7289,g1428,g8992,g579,g6287,g1564,g7351,g1741,g5662,g225,g7309,g281,g7766,g1308,g11627,g611,g9930,g631,g5654,g1217,g9823,g1589,g7359,g1466,g8439,g1571,g7353,g1861,g7815,g1365,g7307,g1448,g11594,g1711,g6335,g1133,g6309,g1333,g11635,g153,g8426,g962,g11404,g766,g6799,g588,g6296,g486,g11331,g471,g11469,g1397,g7322,g580,g6288,g1950,g8288,g756,g755,g635,g5656,g1101,g6814,g549,g11044,g1041,g7788,g105,g11180,g1669,g11036,g1368,g7308,g1531,g7340,g1458,g7327,g572,g10877,g1011,g7805,g33,g10867,g1411,g7331,g1074,g6813,g444,g11259,g1474,g8441,g1080,g6806,g1713,g6336,g333,g5651,g269,g7762,g401,g11266,g1857,g11409,g9,g7336,g664,g8782,g965,g11405,g1400,g7324,g309,g5652,g814,g8077,g231,g7319,g557,g11048,g586,g6294,g869,g875,g1383,g7316,g158,g8425,g627,g5657,g1023,g7799,g259,g7755,g1361,g1206,g1327,g11633,g654,g8067,g293,g7770,g1346,g11656,g1633,g8873,g1753,g5666,g1508,g7329,g1240,g7297,g538,g11326,g416,g11269,g542,g11325,g1681,g11040,g374,g11440,g563,g11050,g1914,g8284,g530,g11328,g575,g11052,g1936,g9355,g55,g7778,g1117,g6299,g1317,g1356,g357,g11509,g386,g11263,g1601,g7363,g553,g11046,g166,g7747,g501,g11334,g262,g7758,g1840,g8694,g70,g7783,g318,g5646,g6818,g794,g6800,g36,g10870,g302,g7773,g342,g11513,g1250,g7299,g1163,g6301,g1810,g2044,g1032,g7800,g1432,g8990,g1053,g7792,g1453,g7326,g363,g11511,g330,g5650,g1157,g6303,g1357,g6330,g35,g10869,g928,g8569,g261,g7757,g516,g11337,g254,g7759,g778,g8076,g861,g4190,g1627,g8871,g1292,g7293,g290,g7769,g1850,g5671,g770,g7288,g1583,g7357,g466,g11468,g1561,g7350,g1527,g4899,g1546,g7345,g287,g7768,g560,g11049,g617,g8780,g17,g4894,g336,g11653,g456,g11466,g305,g5643,g345,g11642,g8,g2613,g1771,g7811,g865,g8275,g255,g7751,g1945,g9356,g1738,g5661,g1478,g8442,g1035,g7787,g1959,g4217,g1690,g6844,g1482,g8443,g1110,g6817,g296,g7771,g1663,g11034,g700,g8431,g1762,g5669,g360,g11510,g192,g6837,g1657,g10875,g722,g9346,g61,g7780,g566,g11051,g1394,g7809,g1089,g6809,g4897,g1071,g6804,g986,g11473,g971,g11470,g6338,g143,g7746,g1814,g9825,g1038,g7797,g1212,g1918,g9353,g782,g8273,g1822,g9826,g237,g7306,g746,g2638,g1062,g7795,g1462,g8438,g178,g7748,g366,g11512,g837,g4184,g599,g9819,g1854,g11408,g944,g11398,g1941,g8287,g170,g8422,g1520,g7334,g686,g9342,g953,g11401,g1958,g6339,g40,g10775,g1765,g3329,g1733,g10882,g1270,g7303,g1610,g6845,g1796,g8280,g1324,g11632,g1540,g7343,g1377,g7312,g4898,g491,g11332,g1849,g5670,g213,g7313,g1781,g7813,g1900,g9351,g1245,g7298,g108,g11593,g630,g7287,g148,g8427,g833,g4183,g1923,g8285,g936,g8571,g1215,g6315,g1314,g11629,g849,g4187,g1336,g11654,g272,g7763,g1806,g8573,g826,g8568,g1065,g7796,g1887,g8281,g37,g10871,g968,g11406,g1845,g5673,g1137,g6310,g1891,g9350,g1255,g7300,g257,g7753,g874,g9821,g591,g9818,g731,g9347,g636,g8781,g1218,g8276,g605,g9820,g79,g7776,g182,g7749,g950,g11400,g1129,g6308,g857,g4189,g448,g11258,g1828,g9827,g1727,g10880,g1592,g7360,g1703,g6843,g1932,g8286,g1624,g8870,g26,g4885,g1068,g6803,g578,g6286,g440,g11260,g476,g11338,g119,g7745,g668,g9340,g139,g8418,g1149,g6305,g34,g10868,g1848,g7366,g263,g7760,g818,g8274,g1747,g5664,g802,g6802,g275,g7764,g1524,g7338,g1577,g7355,g810,g7786,g391,g11264,g658,g9339,g1386,g7318,g253,g7750,g9822,g1125,g6307,g201,g7304,g1280,g7295,g1083,g6807,g650,g8066,g1636,g8874,g853,g4188,g421,g11270,g762,g6798,g956,g11402,g378,g11441,g1756,g5667,g589,g6297,g841,g4185,g1027,g7798,g1003,g7803,g1403,g8991,g1145,g6312,g1107,g6816,g1223,g8277,g406,g11267,g1811,g11185,g1642,g11183,g1047,g7790,g1654,g10874,g197,g6835,g1595,g7361,g1537,g7342,g727,g8434,g999,g7804,g798,g6801,g481,g11324,g754,g4895,g1330,g11634,g845,g4186,g790,g8567,g1512,g8449,g114,g1490,g8445,g1166,g6300,g1056,g7793,g348,g11506,g868,g1260,g7301,g260,g7756,g131,g8420,g7,g2731,g258,g7754,g521,g11330,g1318,g11630,g1872,g9348,g677,g9341,g582,g6290,g1393,g7320,g1549,g7346,g947,g11399,g1834,g9895,g1598,g7362,g1121,g6306,g1321,g11631,g506,g11335,g546,g11043,g1909,g9352,g6298,g1552,g7347,g584,g6292,g1687,g11042,g1586,g7358,g324,g5648,g1141,g6311,g1570,g4900,g1341,g11655,g1710,g4901,g1645,g11184,g115,g7321,g135,g8419,g525,g11329,g581,g6289,g1607,g7365,g321,g5647,g67,g7782,g1275,g11443,g1311,g11628,g1615,g8868,g382,g11442,g1374,g6825,g266,g7761,g1284,g7294,g1380,g7314,g673,g8428,g1853,g5672,g162,g8424,g411,g11268,g431,g11262,g1905,g8283,g1515,g7333,g1630,g8872,g49,g7774,g991,g7802,g1300,g7291,g339,g11505,g256,g7752,g1750,g5665,g585,g6293,g1440,g8988,g1666,g11035,g1528,g7339,g1351,g11657,g1648,g11181,g127,g8421,g1618,g11611,g1235,g7296,g299,g7772,g435,g11261,g64,g7781,g1555,g7348,g995,g7801,g1621,g8869,g1113,g6313,g643,g8064,g1494,g8446,g1567,g7352,g691,g8430,g534,g11327,g1776,g7812,g569,g10876,g1160,g6302,g9824,g1050,g7791,g1,g8078,g511,g11336,g1724,g10879,g12,g7337,g1878,g8695,g73,g7784,I8854,g4500,I9117,I12913,g7845,g11354,I17179,I10891,I10941,g6555,I6979,g2888,g5843,I9458,g2771,I5854,g3537,g3164,g6062,I9699,I9984,g5529,I14382,g8886,g7706,I12335,I13618,g8345,I15181,g9968,g6620,I10573,I12436,g7659,g5193,g4682,g6462,I10394,g8925,I14252,I14519,g9106,g10289,I15691,I14176,g8784,I14185,g8790,I16944,I14675,g9263,g2299,I12607,g7633,g3272,g2450,g2547,g9291,g8892,I6001,g2548,I7048,g2807,g10309,I15733,g7029,I11180,g4440,g4130,I9544,g5024,g10288,I15688,I12274,g7110,I9483,g5050,I12526,I6676,g2759,I8520,g4338,g10571,I16236,I17692,g11596,I17761,g11652,I13469,g8147,I14537,g7956,g7432,g3417,I6624,g4323,I11286,g6551,I8031,g3540,g7675,I12300,g8320,I13344,I12565,g7388,I16644,g10865,I11306,g6731,g1981,I7333,g3729,I13039,g8054,g3982,g3052,g6249,I10006,g9259,I15190,g9974,g11426,I17331,I14958,I13203,I5050,I5641,g5121,g1997,g3629,g3228,g3328,I6501,I12641,g7709,I9171,I10898,g8617,g8465,I15520,g10035,I7396,g4102,I7803,g3820,g3330,I6507,g2991,I6233,I9461,g4940,g2244,I5251,g6192,I9923,I10153,g6085,I9734,I12153,g6874,g4351,I7630,I11677,g7056,g10687,I16356,g4530,I7935,g8516,I13717,g5232,g4640,I13975,g8588,g2078,I8911,g4565,g2340,g7684,g7148,I12409,g7501,I12400,g11546,g11519,I10729,g5935,g5253,g4346,I11662,I7509,g3566,I9427,g4963,g3800,g3292,I15088,g9832,g2907,I6074,I12538,I11143,g6446,g6854,I10920,g11088,I16871,I11575,g8299,I13255,I9046,g4736,g6941,g6503,g2435,I14439,g8969,g4010,g3144,g2082,I6932,g2850,I7662,g3336,I9446,g5052,g5519,g4811,g5740,I9302,I5289,I9514,g5094,I12589,g2482,I5565,I5658,I15497,g10119,g2629,I14242,I11169,g6481,g3213,I6388,I6068,g2227,g11497,I17510,I13791,g8518,I16867,g10913,I10349,g6215,g10260,g10125,I12442,I8473,g4577,I14349,g8958,g6708,I10689,g10668,g10563,I5271,I9191,g5546,I9391,g5013,g6219,g5426,I15250,g9980,I17100,g11221,I14906,g9508,I14976,g7201,I11427,I14083,g8747,g10195,I15559,I8324,g4794,g6031,I9642,g2915,I6094,I13666,g8292,I9695,g5212,I11363,g6595,I11217,g6529,g6431,g6145,g6252,I10015,I10846,I14394,g4372,I7677,g7049,I11228,I6576,g2617,g10525,g10499,g10488,I16101,I10566,g5904,I13478,g8191,g5586,I8996,g8709,g8674,g2214,I9536,g5008,g6176,I9905,g4618,g3829,I15296,g9995,g4143,I7291,I7381,g4078,I9159,g5033,g11339,I17142,g8140,I13017,I16979,I16496,g10707,I12936,I7847,g3435,I9359,g5576,I13400,g2110,I5002,I15338,g10013,g6405,g6133,g8478,I13678,I16111,g10385,g4282,g4013,g11644,I17736,g7604,I12162,g9768,g9432,g4566,g3753,g7098,I11333,g10893,I16641,I4961,g4988,I8358,I10117,g8959,I14326,I13580,g8338,I9016,g4722,I6398,g2335,g8517,I13720,g3348,g2733,I15060,g9696,I15968,g10408,I5332,g8482,g8329,g2002,I10138,g5677,g11060,g10937,I17407,g11417,I12303,g7242,I9096,I15855,g10336,g2824,I5932,g11197,g11112,g4555,I7964,g5691,g5236,g5229,g7539,I11953,g7896,I12678,g8656,I13941,g9887,I15068,I8199,g6974,g6365,I10069,I14415,g8940,g3260,I6428,g11411,I17274,I10852,g6751,g10042,I15253,g10255,g10139,g6073,I9712,g10189,I15545,I4903,g2877,I6025,I11531,g7126,g10679,g10584,g6796,I8900,g4560,I16735,g10855,g1968,g5879,I9498,I10963,g6793,g10270,g10156,g3463,g3256,g7268,I11505,I11734,I11740,g7030,g10188,I15542,I12174,g6939,I12796,g7543,I9138,g7419,g7206,I15503,g10044,I17441,g11445,g6980,I11127,I17206,g11323,g4113,I7255,g6069,I9706,g11503,I17528,g7052,I11235,g8110,g7996,g2556,g4313,g3586,I16196,g10496,I7817,g3399,g8310,I13314,g10460,I15971,g2222,g6907,I13373,g8226,I6818,g2758,I7423,I6867,g2949,I9880,g5405,g10093,I15326,I10484,g6155,g9845,g9679,g3720,I6888,g10267,g10130,g10294,I15704,I11800,g7246,g4908,g4396,g5111,I8499,g11450,I13800,g8500,g5275,g4371,I11417,g6638,I17758,g11647,g3318,g2245,g11315,I17108,g4094,g2744,I17435,g11454,g10065,I15293,I5092,g8002,I12832,g5615,I9043,g4567,g3374,I8259,g4590,g11202,g7728,I12369,I10120,I14312,g8814,I9612,g5149,I16595,I9243,g5245,g11055,g10950,g3393,g9807,g9490,g11111,g10974,g4776,I9935,g5477,g4593,I8004,I11964,g6910,I7441,g3473,I15986,g10417,g3971,I7104,g7070,I11289,g2237,g6399,I10305,g5284,g4376,I11423,g6488,g7470,g6927,I15741,g7897,g7712,g7025,g6400,I6370,g2356,g7425,g7214,I11587,g6828,g2844,I5966,I12553,g7676,I12862,g7638,I8215,g3981,I10813,g6397,g11384,I17209,I14799,g9661,I6821,g3015,g2194,g10160,I15476,I10801,g11067,I14531,I12326,g8928,I14257,g3121,g2462,I16280,g10537,g4160,I7303,g3321,I6484,g2089,I4917,g4933,I8298,I14973,g9733,I5789,I16688,g10800,I11543,g6881,g5420,g4300,I15801,g10282,I12948,g8019,I15956,I12910,g4521,I14805,g9360,I10132,g2557,g4050,I7163,I13117,g7904,I12904,g7985,I4873,g8785,I14090,g4450,g3914,g5794,I9394,g9097,g2071,g7678,I12307,g6144,I9857,I11569,g6821,g3253,I6417,I7743,g3762,g6344,I10251,g3938,I11641,I15196,I14567,g10201,g10175,g7406,I11786,g10277,I15675,g2242,I5245,I9213,g4944,g3909,g2920,I6106,g2116,g7635,I12245,I4869,I13568,g8343,I13747,I15526,g10051,I13782,g10075,I15302,g4724,I10036,I7354,I12463,I5722,g2075,g7682,I13242,g8267,I17500,g11478,g6694,I10663,g4379,g3698,g3519,I12568,I11563,I7411,g4140,g8295,I13239,g2955,I6156,I8136,g4144,g5628,I9062,I6061,g2246,I12183,g7007,g6852,I10914,I11814,g7196,g5515,g4429,I6461,g2261,g5630,I9068,I12397,g7284,g2254,g2814,I5916,I17249,g4289,g4777,g3992,I11807,g11457,I17424,I9090,g5567,g4835,I8192,I14400,g8891,g2350,I5424,I12430,g9267,g9312,I14509,I13639,g8321,g2038,I8943,g4585,I16763,g10890,I12933,g7899,g7226,I11464,g8089,g7934,g10352,I15820,g2438,I11293,g6516,I13230,g8244,g2773,I5858,g4271,I6904,g2820,I12508,g7731,I11638,g6948,I12634,g7727,g10155,I15461,I17613,g11550,g10822,I16534,I4786,I6046,g2218,I9056,g4753,g6951,I11097,g10266,g10129,I8228,g4468,I14005,g8631,g10170,g10118,I8465,g4807,I16660,g10793,g7045,g6435,I10538,g5910,I8934,I5795,g7445,I11845,g6114,I9795,I5737,g2100,I6403,g2337,I5809,I10201,I7713,g3750,g9761,g9454,I11841,I11992,g7058,I11391,g6387,I9851,g2212,I13391,g8178,g6870,I10952,g4674,I8050,g8948,I14299,g3141,g2563,I6391,g2478,I5672,g10207,g5040,I8421,I5077,g1983,I10873,g3710,g3215,g7369,g7273,g7602,I12156,g10167,g10194,g10062,g10589,I16252,I16550,g10726,g4541,I7946,I11146,I17371,g11410,I17234,g11353,g7920,g7516,I11578,g6824,I12574,g7522,g10524,g10458,g2229,I15157,g9931,I16307,g4332,I12205,g6993,I12466,I6159,g2123,g11157,g4680,g6136,I9845,g8150,I7444,g4353,I7636,I10231,g8350,I13430,I13586,g8356,I15365,I8337,g4352,I13612,g6594,I10560,g11066,g4802,g3337,I13442,g8182,g8009,I12849,I5304,I15362,I6016,g2201,I6757,g2732,I12544,I9279,g5314,I9105,I10828,g5875,g5361,g6943,I11079,I16269,g10558,I9720,g5248,I12592,g10616,I16289,g4558,g3880,I9126,I13615,g8333,g7415,I11797,g7227,I11467,I9872,g5557,g10313,I5926,g2172,g8358,I9652,I5754,g2304,I10991,g6759,I15763,g10244,I11275,g6502,g10276,I15672,I17552,I8268,I7760,g3768,I16670,g10797,I11746,g6857,g8241,g10305,I15725,g10254,g10196,g4511,g10900,I16656,g9576,I14713,g2837,g2130,g10466,I15989,g5884,I9505,I5044,g6433,g5839,I9452,g8229,g7826,I6654,g2952,g2620,g1998,I12846,g7685,I5555,I14552,I8815,g4471,g10101,I15335,g10177,I15523,I16667,g10780,I13806,I7220,I5862,g2537,I9598,g5120,I7779,g3774,I17724,g11625,I10907,g7502,I11882,I8154,g3636,I10584,g5864,I17359,g11372,g3545,I6733,I15314,g10007,I17591,I15287,g6195,g3331,g6137,I9848,I9162,g6395,I10293,g3380,g5143,I10234,I16487,g10771,g6913,I11021,g10064,I15290,g11287,g11207,I15085,g9720,g2249,I9625,g4580,I10759,g5803,g11307,I17092,g11076,I16843,I9232,g7188,I11408,g7689,I12322,I17121,g11231,g11580,I11773,I10114,g5768,I9253,I9938,g5478,I16592,g11054,I10831,I9813,g5241,g2344,g5693,I9224,g11243,I17344,g11369,g3507,g3307,g4262,g2298,I5336,g2085,I7665,g3732,g10630,I16311,g11431,g6859,I10937,g7028,g6407,I6982,g2889,I10057,I15269,g9993,g10166,I15494,I11183,I12583,g7546,I9519,g4998,g7430,g7221,I15341,g10019,I5414,I16286,g10540,I7999,g4114,g2854,I5986,I17173,g11293,I5946,g2176,I10849,g6734,g11341,I17146,I7633,g3474,g4889,I8240,g2941,I6118,g6248,I10003,I17767,g9258,g3905,g10892,I16638,I14955,I14561,g3262,I8293,g4779,I10398,g5820,I13475,g8173,I16941,I12627,g3628,g3111,I10024,I7342,g6081,g4977,I10855,I10141,g5683,g4375,g3638,I10804,g6388,I5513,g3630,I6789,g8788,I14097,I11222,g6533,I12282,g7113,I16601,g10806,g5113,I8503,g6692,I10659,I16187,g10492,g6097,I9754,I7732,g3758,g7910,g7460,I12357,g7147,g2219,g9893,I15082,g2640,g1984,g6154,I9875,g4285,g3688,g6354,g5867,g2031,g10907,I16673,g5202,g6960,I11112,I15694,g10234,I5378,g2431,I5510,I15965,g10405,g2252,g2812,g2158,I7240,g7609,I12177,I10135,I11572,g8192,g2958,I6163,g8085,g7932,g10074,I15299,I8462,I13347,g8122,g9026,g8485,g8341,I7369,g5494,g4412,I6941,g2005,g7883,I7043,g2908,g4384,I7707,I9141,g5402,I9860,I8982,g4339,I9341,g10238,g10191,I16169,g10448,I9525,g5001,I14361,g8951,g2829,I5943,g11619,I17675,g2765,g2184,I14964,g11502,I17525,I12439,g2217,I13236,g8245,g7066,g7589,I12099,g4424,g3040,g2135,g4737,g3440,I11351,g6698,I13952,g8451,g5593,I9013,g6112,I9789,I13351,g8214,g6218,I9965,I10060,g3041,I10195,g11618,I17672,g9984,I15184,I11821,g7205,g10176,g10185,g10040,g10675,g10574,I16479,g10767,g10092,I15323,I10048,g5734,I16363,g10599,I16217,g10501,g3323,g2157,I15278,g10033,g7571,I12035,I11743,g4077,I7202,g6001,g7048,I11225,g10154,I15458,g2270,I5311,I5798,I17240,g11395,g7711,I12344,g4523,g3546,I10221,g6117,I11790,g8520,I13729,I17444,g8219,g2225,I5210,g8640,g8512,g10935,g10827,I5731,g2073,I4879,g2796,g2276,I16778,I6851,g2937,I7432,I7697,g3743,I10613,g6000,I11873,g6863,g10883,g10809,I17755,g11646,I11647,I7210,g2798,I12487,g5521,g3528,I14323,I16580,g10826,I17770,g11649,I16775,I8429,g2124,g3351,I6535,g5641,I9084,I17563,g11492,g2980,g6727,g5997,g8376,I5632,I5095,I6260,g2025,g2069,I9111,g5596,I11420,g4551,g3946,I15601,g10173,I9311,g4915,I15187,I12248,I13209,g8198,g4499,I8848,g4490,g2540,I5655,g7538,I11950,I13834,g8488,I5579,I12505,g5724,I9268,g9027,I14418,g2206,I5171,I12779,g7608,g10729,g6703,I10678,I9174,g4903,I5719,g2072,g10577,g10526,g11648,g7509,I11889,g9427,g9079,I10033,I7820,g3811,g4754,I16531,g10720,g10439,g10334,g6398,I12081,g6934,g5878,g5309,I11058,g7662,I12279,g4273,I16178,g10490,I12786,g7622,I17633,g11578,I9135,g5777,I9365,I10795,g6123,I13726,g8375,g7467,g1990,g2248,g8225,I17191,I17719,g11623,I11614,g6838,g8610,g8483,I6367,g2045,I9180,g4905,I12647,I16676,g10798,I16685,g10785,I11436,I9380,g10349,I15811,I14540,I16953,g11082,I13436,g8187,I9591,g5095,I16373,g10593,g4444,I7800,g8473,I13669,g2199,I17271,g2399,g9763,g7093,I11326,I12999,g7844,g3372,I10514,I12380,g7204,g10906,I15479,g10091,I13320,g8096,g10083,I15311,I9020,g4773,g8124,g8011,g10284,g7256,I11489,I12613,g8324,I13354,g11479,I17470,I6193,g2155,I11593,g6830,g3143,I6363,g11363,I17188,g3343,g2779,I11122,g6450,g2797,g2524,I13122,g7966,I6549,g2838,g4543,I10421,g5826,g6443,I6738,I6971,g2882,g6716,g5949,I14421,g8944,I5254,g6149,I9866,g3988,I6686,g6349,I10258,g7847,I12638,g3693,I11034,g6629,I10012,g5543,g3334,I6517,I5725,g2079,g7197,I9617,I15580,I13797,I6598,g2623,g7021,I11162,g4729,g4961,I8333,g7421,I15415,I5410,I8211,g5300,I10302,I10541,I6121,g2121,g1963,g110,I17324,g11347,g7263,I11498,I14473,g8921,g2207,I5174,g10138,I15412,I17701,g11617,I10789,I12448,g7530,I13409,g8141,I17534,g11495,g3792,I7017,g5353,I8820,g8849,g8745,g2259,I5292,g6241,I9992,g2819,g2159,I11635,g6947,I10724,g6096,g11084,I16863,g4414,I7752,I10325,g6003,g11110,g3621,I6754,I6938,I7668,g3733,g2852,I5982,I7840,g3431,I16543,g10747,g10852,g10740,I14080,I8614,g6733,I10535,I12026,g7119,I10434,I16938,g2701,g2040,g3113,I6343,g7562,g6984,I14358,g8950,I7390,g4087,I10946,g6548,g8797,I14116,g6644,I10601,g4513,g7631,I12235,g7723,I12354,g6119,I9810,I9973,g5502,I12616,g5901,I4920,g8291,I13227,g11373,I17198,g3094,I6302,I7351,g4436,I10864,g4679,I17764,g4378,g7605,I12165,g5511,g6823,g3518,I10682,g6051,g10576,I9040,g8144,I13027,g8344,I13412,g6717,I10706,I9440,g5078,I17302,I13711,g8342,I16814,g10910,I12433,g7657,g4335,I7612,I9123,g4890,I11109,g6464,I12418,I7363,I9323,g5620,I13109,g7981,g4288,I11537,g7144,g4382,I16772,g10887,g3776,g2579,g6893,g5574,g10200,g10169,g2825,I5935,g2650,g2006,g10608,I16283,g10115,I15353,g6386,I10282,g7585,I17447,I5684,I8061,g3381,g4805,g2643,I5963,g2179,I7810,g3799,g7041,g6427,g4005,g10863,g2008,I13606,g8311,I12971,g8039,I11303,g6526,I10081,g3663,g6426,I10340,g11423,g2336,I16416,g10664,g7189,g5278,I7453,g3708,g6170,I14506,g8923,g7673,I12296,I9655,g5173,g6125,I9822,I5707,g2418,I14228,g3521,I14306,I16510,g10712,g5262,g3050,I11091,g6657,g10973,I16720,g5736,I9296,g6382,I10099,I11071,g7669,I12286,I17246,g11543,g3996,g10184,g10039,I12412,g7520,I8403,g4264,g10674,g8314,I13326,g5623,I9053,I12481,I7157,I11255,I12133,I5957,g2178,I7357,g2122,g2228,g7531,I11929,g4095,I7233,g9554,I14697,I14182,g2322,I10927,g6755,g7458,g7123,g5889,I12229,I6962,g2791,g4495,I7886,I9839,g5226,g2230,g4437,g3345,I7244,g11514,g7890,g7479,g8650,I13933,I13840,I16586,g10850,g3379,I15568,g10094,g10934,g6106,I9773,g5175,I10177,g7505,g3878,g11242,I5098,g8008,I10240,g5937,g7011,g4719,g10692,I9114,I6587,I10648,g6030,I15814,g10202,g8336,I13388,I14903,g9507,I5833,g2103,g6121,g5285,g4355,g6461,I10391,I15807,I15974,g10411,I8858,g4506,g2550,g7074,I11299,g10854,g3271,I6443,g10400,g10348,g2845,g2168,I9282,g5633,I15639,g10179,I10563,g6043,I5584,g10214,I15586,g9324,I14970,g2195,g4265,g3664,g10001,I9988,g5526,I10343,g7697,g2395,g2891,I6055,g5184,I5395,I11483,g6567,g2913,I6088,g10329,I15775,g10186,g4442,I6985,g2890,g6904,I11008,g6200,g11638,g10539,I16184,g4786,g6046,I9669,I7022,I8315,g4788,I8811,g4465,I10370,I12981,I7118,g8289,g9529,I14672,g4164,I7311,g10538,I16181,g4233,g5424,I8865,I14549,g6660,I13949,g6403,g6128,g8203,I9804,g5417,g2859,I5995,g3997,I7131,I15510,I14570,I9792,g5403,I6832,g2909,g4454,g8033,I12875,I17549,g6191,g5446,g7569,I12029,I9177,g4296,I7559,I11904,g6902,I10633,g6015,g6735,g5231,I17318,g11340,g3332,I6513,I11252,g6542,g10241,g10192,g9260,g6695,I10666,I10719,I13621,g8315,g3353,I7735,g3759,g2808,I14191,g8795,I12953,I17616,g2342,I5406,I7782,g3775,g6107,I9776,I17540,g11498,I12857,g11014,I10180,g3744,g6536,I10456,I4883,g5205,g4366,g10159,I8880,g4537,g2255,I5276,I5728,g2084,g7688,I12793,g7619,g2481,I9202,g8195,g7976,I12776,g8137,I13010,I14239,g8337,g10235,g4012,I7154,g6507,I16193,g10485,I17377,g2097,I4935,I12765,g10683,g10612,g5742,I9308,g2726,g2021,I7746,I11397,g6713,I13397,g8138,g2154,I5067,g6016,I9632,I12690,g7555,I7384,I5070,g2960,I6173,I10861,g5980,I9567,g5556,g8807,I14140,I14573,g9029,I8237,I11367,g8505,g11412,I11626,I10045,g5727,g6115,I9798,g6251,I7330,I10204,I10843,I15275,g9994,I7674,I14045,g8603,I17739,g11641,g4787,g3423,g4728,I16784,I16616,g5754,I9332,g5800,I16475,g10765,g6447,g6166,I10388,g5830,I8234,g4232,I12445,I14388,g8924,I8328,g4801,g11305,g10972,g3092,g2181,I14701,g6126,I14534,g9290,g4281,g5493,g5613,g4840,I10958,g8142,I13023,g2112,I13406,I15983,g10414,g2267,I17698,g11616,I16766,g8255,g7986,g8081,g8000,g8481,g2001,g7924,g7220,I11456,g5572,I8989,g5862,I9479,I12502,I4780,I6040,g2216,g10522,I15517,I13574,g8360,g2329,I5383,g8354,g8717,g7023,I11166,I7952,g10206,g10178,I5801,I7276,g2861,g9670,I16781,g4791,I8161,g7977,g2828,I5940,I10075,g10535,I6432,g2727,g2022,g3736,I6924,g5534,g4545,g5729,I11731,g10114,I15350,I16175,g9813,I14948,I15193,g6417,I13051,g8060,g9987,g6935,I11065,g11193,g7051,I11232,g10107,I11756,g7191,g2221,I5198,g3076,I6282,I13592,g8362,g8783,g8746,g10058,I11629,I12232,g7072,I6528,g3274,I16264,g10557,I16790,I8490,g4526,I7420,I6648,g2635,g8218,I9658,g5150,g8312,I7546,g4105,I9829,g5885,g10345,g7999,I12825,g7146,I5445,I11686,I10162,g5943,I12239,g4049,g3375,I6569,g8001,I12829,I12261,g7078,g4449,g3722,I6894,I8456,g4472,g7103,I11338,g5903,g4575,g10848,I16546,g11475,I17466,g8293,I13233,g8129,g8015,I6010,g2256,g2068,I4866,I11152,g6469,I13367,g10141,I15421,g7696,g10804,I16514,I10810,g4098,g3500,I6690,I15437,g10050,I16209,g10452,I8851,g4498,g8828,g8744,g11437,I17362,g2677,g2034,g10263,g10127,I12424,I9981,g5514,g8727,g8592,g5679,I9194,g7508,g6950,g3384,g10332,I15782,g6213,I13837,g7944,g7410,I15347,g10135,I15403,g7521,I17164,I8253,I7906,g3907,g2349,I5421,g7043,I11214,I12499,g7725,I11405,g6627,g5288,g4438,I14528,g3424,g2896,I9132,g4893,g10361,g10268,g3737,g2834,g7443,g4935,g9525,g9257,I9153,g5027,I9680,g5194,I10147,g5697,I10355,g7116,g5805,I9409,g5916,I9550,I11596,g2198,g2231,g4268,I7523,I7771,g3418,I16607,g10787,g2855,I5989,g4362,I7651,g6901,I14355,I12989,g8043,g11351,I17170,g3077,g2213,g5422,g4470,g7034,I11191,I10825,g6588,g4419,I7763,I9744,g5263,I12056,g6929,g5857,I9893,g8624,g8486,g3523,g2971,I14370,g8954,g8953,I10858,g6688,I13020,g8049,I13583,g4452,g3365,I8872,g4529,I15063,g9699,g2241,I11394,g6056,g5947,I9585,I11689,g11063,I11046,g6635,I10996,g6786,I12271,g7218,g7681,g6649,I10610,g4746,g8677,I13962,I10367,g6234,g5824,I9901,g7101,I14367,g8884,g10864,g3742,I6929,g7914,g7651,g8576,I13819,g7210,I11440,I8080,I16292,g10551,g2644,I10671,g4730,g8716,I17546,g11500,g8149,I13036,g10947,I16708,g4504,I7899,I11357,g6964,g6509,I13427,g2119,I5031,I10039,g5037,I8414,I13357,g8125,I12199,g7278,I7372,g3226,g9311,g11422,I17321,g7035,I13105,g7929,I9120,g4385,I7710,g7413,g5102,I8476,g2258,I14319,g8816,g2352,I5430,g2818,I5922,I7140,g2641,g6063,I12529,g2175,g2867,I6007,I16635,g10862,I15980,g11208,g11077,I7843,I13131,I8256,I14040,I7478,g5719,I9259,g4425,I12843,g7683,I16717,I15235,I5388,I7435,g3459,g7936,g11542,g11453,I17416,g5752,I9326,I13803,g8476,g3044,I6256,g2211,g9310,I10096,g2186,I11599,g6720,I10713,g4637,g6118,I9807,g3983,g3222,g11614,I17662,g7601,g5265,g11436,g3862,g5042,I15320,I14989,g6652,g4678,g6057,I10901,I15530,g11073,g4331,I7606,g3543,g3101,g2170,g2614,g1994,I12490,g7922,I12712,g2125,I5053,g8319,I13341,g11346,I17161,I15565,g2821,I5929,g9268,I15464,I6965,g2880,g4766,g7033,I10739,g5942,I7249,g8152,I13043,g10421,g10331,I16537,g10721,g4305,g6971,g6517,g8051,I12258,I6907,I6264,g2118,I16108,g10383,g6686,I10651,g10163,I15485,I14010,g7597,g5296,I11249,g6541,I5638,I14645,g9088,g2083,I6360,g4748,I16492,g10773,I13482,g8193,I5308,g97,I11710,g7020,I12517,I4992,g4755,g10541,I16190,I10698,g5856,I9816,I15409,I7002,g8186,g10473,g10380,g4226,I11204,g6523,g6670,I7402,g4121,I17268,I6996,g2904,I7099,I13779,g8514,I7236,g3219,I15635,I16982,g8599,g8546,g7995,I12817,g2790,I17265,g7079,I11312,I11778,g3903,I7070,g5012,I8388,g9100,I13194,I10427,g4445,I10018,g2061,g2187,g6938,I11068,I7336,g4373,I7680,I16796,g11016,I16172,g4491,I12986,g7190,I11412,g8325,g6925,g7390,g6847,I12878,g5888,I13945,I12171,g6885,g10121,I15371,I14373,g3436,g4369,I13212,I7556,g4080,g4602,I8011,I11879,I17450,g3378,I6572,g5787,I9383,I9424,g5404,I17315,g11393,g10344,I15798,I9737,g5258,I6065,g2200,g6552,g5733,I11716,g2046,I17707,g4920,I5827,g2271,g2446,g4459,I17202,g11322,g3335,I6520,g8265,g8332,g4767,I8123,I7064,g2984,g11575,g11561,g2003,g5281,g4428,g3382,I6580,I9077,g4765,g4535,I6611,g2626,I8506,g4334,g2345,g10120,I17070,g11233,g8106,g7950,g11109,g8306,I13290,g2763,I5847,g2191,g2391,I5478,g6586,I12919,g8003,I6799,g2750,I11932,g6908,g3749,I14101,I9205,g11108,g2695,g2039,g9666,I14793,I12901,g5684,I8275,I8311,g4415,g5639,I9080,I14127,g8768,I17384,I12595,I11737,g10134,I15400,I7295,I11961,g7053,I16553,g10754,g5109,I8495,g5791,g3798,I13448,I9099,I5080,I11824,I14490,g8885,g6141,I9854,g8622,g6570,g6860,g6475,I11238,g6585,I14558,I5662,g9875,I15036,I13595,g9530,g6710,I10693,g5808,g5320,I5418,g2858,I5992,I12598,g7628,I7194,I14376,I14385,g8890,I7426,I8985,g4733,g11381,g4721,g2016,g2757,I5837,I13636,g7568,g5759,g5271,I10888,g6333,I6802,g2751,g3632,g3095,g3037,I12835,I14888,g10515,g3437,g7692,I9273,g5091,g6045,I17695,g3102,I4924,g3208,I6381,g7912,g8145,I13030,I13415,g2251,g2642,g1988,I12159,g7243,I11719,g2047,I12532,g7594,g7984,I13114,g10927,g9884,g6158,I9883,g3719,I12783,g7590,g11390,I17219,I13723,g8359,g5865,I9486,I13978,g2275,I6901,I11149,g6468,g2874,I6022,g7519,g3752,I6947,g10782,I11433,g6424,I16847,g10886,I11387,g6672,g5604,I9032,I13433,g8181,g5098,g2654,g2012,I11620,g6840,g5498,I8919,g5230,g6587,g5827,g4388,I7719,g10491,g10903,g6748,I13457,g6111,I9786,I10084,I10192,I7465,g10604,g8858,g8743,g4671,g3354,I6028,I7776,I5646,I10546,g5914,g5896,g4430,I14546,I7438,g3461,g3364,I7009,g5700,I8204,g3976,I12631,g7705,g8115,g7953,g4564,g8251,I13166,I13329,g10025,g2017,I10111,g2243,I5248,g3186,g3770,g6239,g10794,I15536,g10111,g10395,g10320,g5419,g9804,I14939,g10262,g10142,g10899,g10803,g6591,I10553,g6411,g4394,I5101,I14194,g3532,g2234,g6853,I10917,I10126,g5682,g6038,I16574,g10821,g4638,g2328,I12289,g7142,I6968,g2881,g6420,I10334,g11621,I17681,I5057,I15551,g2542,I8973,g4488,g2330,g7735,I12384,g4308,g3863,g6471,I17231,g11303,I12511,g6559,g5758,I12571,g3012,I6247,I11011,g6340,I5751,g2296,g8595,g6931,I11055,g5728,I9276,g5486,g4395,I10296,g6242,g7026,g5730,g5504,g7949,g7422,I7468,I16950,g3990,g2554,g4758,g4066,I7191,I13188,g10781,g4589,I7996,g5185,g5881,g7627,I12223,g9094,I5041,g5198,g4466,I7833,g1992,g6905,I5441,g3371,g11062,g7998,I12822,g10247,g4165,g4365,I13627,g8326,g5425,g10389,g10307,g10926,g6685,I13959,I13379,g8133,I17543,g4711,g6100,I9759,g6445,I17716,I10159,g7603,g4055,g7039,I9749,g5266,g10388,I8351,g8234,g2902,g7439,I11833,g8128,I12993,I13364,g7850,g10534,g10098,I15332,I17456,g4333,I7837,g4158,g8330,I13370,g10251,g10272,g10168,g2090,g4774,I7462,g3721,g5415,I13096,g7925,g2166,g6750,g9264,I14477,I6424,g7702,I7405,g5678,I10503,g5858,I16413,g10663,g10462,I15977,g3138,I6356,g8800,I14123,I14503,g8920,I8410,g4283,g2056,I4859,I16691,g10788,I14579,g3109,g3791,I7014,g2456,g7919,g7512,g10032,I15232,g2529,g2649,g10140,I15418,g4780,I8839,g4484,g6040,g2348,I6077,g11574,g11452,I17413,I16802,I9199,g5766,I9346,I8487,g4509,g6440,g6150,g1976,g11205,I6477,g7952,g7427,g9450,g5305,g5801,I5734,I6523,I4820,I17243,g11396,I5435,g2851,I5979,g2833,I12559,g7477,I14315,g8815,I6643,g3008,g8213,I10819,g6706,g11311,I10910,I9102,I9208,g5047,g3707,I14910,g9532,g7616,I12196,g7561,I12015,g4067,I6958,I8278,g8805,g5748,I9320,I10979,g6565,g2964,g4418,I9869,g4467,I15072,g9713,I14979,g9671,g4290,I14055,I16583,g7004,g11072,I17773,g11650,I15592,I15756,g7527,I6742,g3326,g4093,g2965,I8282,g4770,g6151,I12457,g4256,g6648,I10607,g9777,g9474,I11970,I10384,g5842,g10162,I15482,g3715,I9265,g5085,I16787,g10896,g11350,I5713,g2436,g10204,g8056,g7671,I13317,g8093,I12610,I7360,g2906,g8529,I13738,I14094,g8700,g4381,g7476,g5396,g8348,I13424,I12255,g7203,I6273,g2872,I16105,g10382,g10629,g10583,I10150,g5705,g5169,g4596,I7408,g8155,I13048,I13002,g8045,g8355,I13445,g10220,g5007,I8379,I13057,g7843,g2652,g2057,g7376,I13128,g2843,g10911,I11608,g2989,g3539,g4263,I13245,g8269,g7042,I16769,g10894,g5718,I9256,I12460,I12939,g5767,I9349,g10233,I13323,I7176,I5976,g2549,g2853,I10526,g6161,I12907,I5952,g6172,I10093,g7617,g3861,g7906,I12694,I17258,g5261,g10591,I16258,I6543,g3362,I6546,g3419,g3104,I7829,g3425,g6667,I10630,g4562,I7973,g6343,I10248,I16439,I14564,g10355,I15829,I10105,I12478,g6566,g7027,g4631,g10825,g6732,I15583,g10157,g9802,g1999,g6537,g4257,g6134,I13338,I14188,g5221,g2232,I5221,g10172,I16799,g3086,g5203,g2253,g3728,g2813,I5913,I9029,g4781,I14077,g8758,g4902,g6080,I9371,g5075,I10822,I15787,g10269,I6414,g3730,I6080,I9956,g5485,g6059,g3385,g11357,I17182,g7991,I12809,g10319,g4441,g6113,I10198,I11309,I11668,I10102,g10891,I13831,g8560,g10318,I15752,g4089,I5588,g8121,I12978,g10227,g7907,g7664,I6436,g2351,I6679,g4673,g6202,g8670,g8551,g5689,I9216,g4757,I9684,I11194,I15768,g10249,g5210,I9639,g5126,g7959,I12751,I10066,g5778,I9338,g8625,g8487,g7082,I11315,g2586,g1972,g5216,I17410,g11419,g6094,g6578,I16647,g10866,I15281,g10597,g4669,I8724,I10495,g4368,I11989,g6919,I17666,g11603,I10885,g6332,g4231,I6510,g10203,I14876,g9526,I11611,g7656,I12265,g4772,g3406,I11722,I7399,I15263,g3635,I6812,g4458,g2570,g2860,I5998,g2341,I5403,g9262,g3682,g6593,I10557,g5344,g8519,g3105,g7915,g7473,g3305,I6474,g10281,g98,I4783,g2645,g1991,I8835,g7677,g10902,g8606,I11450,I15368,g4011,I7151,g9076,g5741,I9305,g3748,g4411,g4734,I11342,g9889,I11345,I10051,I6560,g3212,I8611,g5844,g5638,g6933,I11061,g7663,I11650,g10699,I16376,I12853,I16897,I5240,g2962,I6183,g6521,I10437,I17084,g11249,g4474,g10290,g6050,I9677,g6641,I10598,I11198,g5081,g10698,g2506,I10378,I6037,g2560,g11348,g5883,I10314,g7402,I6495,g2076,I9833,g5197,I11528,I6102,g2240,g10779,I17531,g11488,I7694,I11330,g6571,g3373,I6565,I15778,I12451,g3491,g2669,g2903,I5116,g11081,I16856,I7852,g3438,I7923,g3394,g5066,I8436,g5589,I9001,g6724,I13403,I10054,I9539,g5354,I9896,g5295,g4713,I10243,g5918,I11132,g6451,I11869,g6894,g7877,I7701,g3513,g3369,I6557,I6240,I14522,I15356,I12268,g6878,I10966,I15826,g10205,I6917,g2832,I15380,I4894,g2174,I6661,g9024,I14409,g2374,g7534,g5035,g7556,I16723,g10851,g3767,I6976,g10547,I16206,g9424,g10895,g4076,I9362,g2985,I6217,g9809,I14944,I9443,g6882,I10974,g7928,I10156,I10655,g6036,g10132,g3582,I16387,I17334,g11360,I10072,g6534,g10226,I15598,I16947,g11651,g7064,I11269,g2239,g9672,I13708,g5774,I12683,g3793,g2593,g7464,I11858,I12053,g6928,I13454,g7686,I12520,I16811,g10908,I16214,g3415,g3227,I6406,I7825,g3414,I10807,g2171,I11043,g6412,I6454,g2368,g8055,I17216,g11291,g2420,g6674,I10639,I17558,g7259,I15383,g3209,I13197,g2507,g3246,I15448,g10056,g5509,g4739,g4326,I14694,g4125,g7237,I11477,I9185,I6891,I11602,g6833,I11810,I17255,g6132,I9147,I6553,I4850,g11499,I13068,g6680,I10643,g6209,g5994,g10889,I16629,I16850,g10905,g6918,g7394,g6197,g10354,g2905,g7089,I11322,I12376,g10888,I16626,I10816,g8239,I7366,g9273,g4608,g3726,I12762,I4948,I10278,g5815,g3940,g6558,I12009,g6915,I8262,g4636,I11967,g6911,g8020,I10286,g6237,I5060,g10931,g3388,I6590,g8812,I11459,g11433,I17350,g9572,I14709,g5685,I9237,g8794,I14109,g5397,I5818,I8889,g4553,g11620,I17678,g10190,I15548,g4361,I7648,I9766,g5348,g3428,I6639,I7096,I12454,g7544,I9087,g4970,I9801,g5416,g3430,g7441,I17742,g4051,I7166,g5996,g8047,g11343,I17152,I13918,I16379,g10598,g4127,g4451,g4327,I7600,g11352,I11698,g6574,g2196,g10546,I16203,g7038,I11201,I11444,g6653,g11420,g10211,g9534,I14687,I15162,g6714,g7438,g7232,I12484,g6832,g7009,I17194,I5047,g2632,I7625,g8515,I13714,g10088,I15317,I8285,g4771,g7073,I5840,g2432,g9990,g11481,I16742,g10857,g8100,g7947,g11079,g3910,I13086,I12472,I8139,g3681,g7212,g5723,I14884,I17277,I11817,I10168,g5982,g5817,g7918,g5301,g7967,I15229,I5427,I11159,g6478,g10700,I5765,I9491,g5072,g10126,I8024,g4117,I11901,g6897,g2530,g6736,I13125,g7975,g8750,g6042,g4508,g10250,g10136,g2655,g2013,g4240,I11783,I16793,I9602,I5704,g7993,I12813,g6076,I9717,I4906,I11656,g7122,I6049,g5751,I6955,g3066,I8231,g4170,g4443,g3359,g10296,I15708,I11680,I14340,I17116,g11229,g2410,g9452,I7726,g6175,g4116,I7260,g6871,g2884,g2839,I7054,I6498,I17746,g11643,g3055,I15959,g10402,g7921,g7463,g10197,g4347,I8551,g4342,g3333,I9415,I17237,g11394,g4681,g4330,I12577,g7532,g8151,g8036,g10527,I6999,g8351,I17340,g11366,g4533,I7938,g7848,g8221,I15386,g6184,I9915,g2235,g2343,I9168,I10531,g6169,I17684,g11609,I14179,I7447,I7112,g11301,g11096,I16879,g7620,I12208,I8007,g3538,I6726,I6019,g6140,g10859,I10186,g6110,g6737,I16571,g2334,I10837,I10685,g6054,g5743,g4413,I7749,g5890,g6508,I6052,g2220,I5667,g8956,g6531,g8050,I14224,I16298,g10553,I13224,g8261,g6077,g11429,g5011,I8385,g3067,I13571,g10315,g10243,I9290,g10819,I16525,g11428,I17337,I16682,g3290,g11376,g10171,g10257,g4317,I7586,I13206,I4876,g3093,I6299,g5474,g7192,g6742,g5992,I9608,g7085,I11318,g3763,g6634,I10589,I9188,I10762,g6127,g8667,g3816,g8143,g8029,I13816,g8559,I6504,g3214,I9388,g8235,g11548,g6104,I9769,g9762,g10590,I16255,I6385,g2260,I10171,g10909,g6499,I16261,g10556,g2202,g11504,g4775,I11752,g7032,g8134,I13005,g7941,g8334,I13382,g9265,g2094,I12415,g11317,I17112,I15329,g3397,g8548,g8390,g2518,g4060,g4460,I9564,g3697,I10078,I8885,g4548,g8804,I14133,I14543,g4293,g10150,I16507,I9826,g5390,g7708,I12339,g8294,g10735,g11057,I11898,g8792,I14105,I17347,g3735,g6044,I9665,g1973,g7031,g6413,I8903,g4561,g6444,g11245,g7431,I12601,g11626,g9770,I15562,g6569,g10695,I16366,g5688,I17124,I13489,g8233,I6196,g2339,I5475,I7716,g3751,g6572,g6862,I5949,g7580,g8787,I9108,g10253,g8200,g4479,I7858,I14681,g6712,g5984,I8036,g4294,I10123,g5676,g6543,g4462,g9553,g8767,g3723,g3071,g7286,I11534,I7387,g2197,g4390,g6396,I15962,g3817,g7911,g6563,g8094,g7987,g2050,g1987,I8831,g4480,I17516,g11483,I16432,g10702,g4501,g6729,g6961,I11115,I13794,g5863,g4156,I11713,g7733,I5850,g2273,g7270,I11515,I11049,I6944,I9165,I16461,I9571,g5392,g7610,I12180,g4942,I8308,I14424,g6014,I11296,I12799,g9429,g9082,g22,I4777,g5838,g11289,I10623,g6547,g10256,I17555,g8270,I14391,I16650,g10776,I6373,g2024,I6091,g5183,g7124,g7980,g10280,g6903,I11005,g2777,I5919,I11188,g6513,g7069,I12805,g8171,g5779,g9272,g4954,g4250,g4163,I7308,I6034,g7540,I11956,g8160,g4363,I7654,I16528,g10732,I7577,g4124,I13460,g10898,g5423,I17453,g11451,I11383,g6385,g7377,I11759,I15467,I9647,I5561,g8052,g4453,I13648,g6178,I6767,g2914,g4325,g3368,g9745,g2826,g2799,I17513,g6135,I9842,I9156,g9109,I14452,I10228,g9309,g3531,I8869,g4421,g5127,I8535,g3458,g6182,g11389,I9662,g5319,g8179,g7849,I12644,I16598,g10885,g11056,g8379,I13485,g4912,g8766,g2997,I17657,g7537,g2541,g11080,I16853,g5146,g10708,g3505,I6694,I5970,g2185,g6749,I10756,g2238,I5237,g11432,g3411,I6616,I9093,g7900,g10555,g2209,I12556,I8265,g5696,I9229,I11085,I7984,I5224,I7280,I10237,g6120,I8442,g4464,g7658,I13185,g2802,g11342,I17149,g6205,I5120,g9449,g6560,g8820,g5753,I9329,I8164,I15736,g10258,g10456,g5508,I8929,g11199,I14684,g9124,I17752,I11617,g6839,I13915,g5472,I14364,I9421,g5063,g2162,g5043,g6522,g10314,I15744,I11494,g5443,g6208,I9953,I7790,g3782,g10936,I10165,I15729,I7061,g6579,g5116,g6869,I10949,g7852,g7923,g11320,g4083,g10596,g8339,g8132,g6719,I10710,I13376,I11623,g6841,g7387,g8680,I13965,g10431,g10328,I11037,g8353,I13439,I14130,g8769,I10362,g6224,g2864,g5948,g6917,I11029,I8247,g2208,g8802,I6671,g7886,g4735,I17327,g11349,I7109,g4782,I11155,g6470,I17537,I13418,I13822,g6442,I11590,I8631,g11225,I7345,I16458,g10734,I9605,g4475,g6164,g3769,g2646,g5755,g10335,g7650,I15244,g10031,g4292,g10930,g6454,g11244,I7931,g6515,g3760,g3003,g7008,I13589,g8361,I17381,I7536,I4886,g10131,I15395,I11524,g11069,g4084,g3119,I11836,g4603,g5936,g8600,g8475,g9710,I12469,g4439,I7793,g5117,g6553,I10477,g8714,g11068,g3631,I12120,g10487,I16098,g7972,I12770,I11119,g9025,I14412,g2871,I6013,g10619,I12759,I7757,I16817,g10912,I9673,g5182,I14236,g6556,g3220,I8109,g3622,g2651,g2007,g2302,g4583,I10322,I17390,g11430,g10279,g10158,g7065,I11272,I7315,g6389,I10289,I7642,g7887,g7693,I15792,I9368,g4919,I8290,I10063,g6990,g3694,g10278,g10182,g3977,I6861,g2942,g6888,I10984,g10791,I9531,g5004,g6171,I16295,g10552,g3161,I11704,g7632,g2569,I17522,g11485,I5399,g6331,g6956,I11106,g5597,I9023,I14873,I13809,g8480,I6133,g3051,g2165,I12930,g10069,I13466,g5088,I13674,g2424,I8449,g4469,I12652,g9766,g2809,I5909,g5784,g4004,g5257,g8053,g4518,g7550,I11560,g7037,g10187,I15539,I5824,g2502,I10834,g6715,g3633,I15079,I8098,g3583,g2077,I5218,g7195,g11545,g11444,g7395,I13642,g8378,I11659,g3103,I9074,g4764,g7913,I6538,g2827,g2523,I7272,g1989,g10143,I15427,g11078,I10021,g5692,g5840,I13695,g11598,I17642,g3068,g6109,I12406,g11086,I12586,I7417,I6914,I17252,g8184,g10884,I15817,g10199,I9863,g8139,g8025,g2742,g3944,I15500,g5763,g6707,I13630,I5348,g9091,g4320,g11159,I10274,g5811,g6480,I11665,g3761,I5064,I14112,g10217,I15589,g4277,g6201,I11674,g6795,g6957,g2754,I5830,g4789,g10486,I16095,I17176,I15823,g6449,g8194,g8477,g8317,g6575,g7525,g8523,I13732,g2257,g9767,I14914,g7097,I9688,g5201,g7726,I12363,g5269,g8183,I5740,g7497,g9535,I14690,I10702,g10580,g10530,g2444,g5032,g2269,g10223,I15595,I7213,g9261,I6421,g2346,g4299,g8938,g7579,I6856,g8099,g7990,g4238,I14136,g8775,g8304,I13280,g4891,g8266,g10110,I15344,g2543,g6584,g11017,g6539,I10461,g6896,g5568,g10321,I15759,I5089,I17213,g11290,I12514,g10041,g10531,g10471,g7979,g3413,g5912,I11584,g4738,I11519,I11176,g6501,g7001,I11140,I13191,g10676,g10570,g6419,I10331,g6334,I7456,g3716,g1993,I7284,g6052,g11309,I17096,I7205,g8613,g8484,g10719,I7348,g4056,g6452,I15308,g4478,g2014,g2885,I6043,I9779,g5391,g2946,g4435,g4727,g4082,I12421,g7634,I8406,g4274,g8765,I12366,g3433,g9308,I10108,g6086,g8712,I12012,g6916,I9588,g5114,I12403,I5438,g11377,I14303,g8811,I10971,I12541,g7703,g5174,g10264,I5525,I15374,g9028,g8729,g8961,I14330,I4900,I11501,g6581,I16610,g10792,I14802,g11308,g3060,g8290,I13577,I10381,g5847,I7459,g10554,I14982,g6425,I11728,g7010,I17733,I16679,g10784,I5391,g2979,g4310,g2382,I7318,g3266,g7680,I16124,g10396,I12535,I10174,I15669,g10543,g3784,g11425,g5894,g10117,I15359,g8660,g8946,I14295,g2916,I6097,g5735,I9293,I15392,g10104,g2749,I5815,g3995,g3937,I7086,I10840,g9741,g4002,I7393,g4096,I6531,I11348,g7062,I13083,g3479,g11195,I17482,g6131,g5548,I9144,g8513,I15488,g10116,I15424,g10080,g6406,g10242,I15632,g5475,I8892,g4762,I8116,g2449,I11695,g11424,I9240,g5069,I10592,I11566,g6820,I16739,g9108,I14449,g3390,I14499,g5627,g5292,g9883,g3501,g4340,g5998,I9620,I13385,g2873,I10753,g2095,I11653,g6954,g2037,I13099,g4222,g5603,g2297,g5039,I8418,I4951,g10293,I15701,g2653,g2011,g6922,g5850,g6226,g3704,g10265,g1969,g8357,g6747,g11391,g2719,g2043,g9448,I7909,g3387,g2108,g8818,g4785,g10391,I6480,g5702,g2752,g8649,g9555,g6091,g6071,g3810,g3363,I10904,g8798,I14119,I11354,I11605,g3432,g10579,g10528,g4563,g9774,g4166,I13773,I16277,g10536,g2042,g4295,g10578,g4237,I10317,g6868,g5616,g10783,g8632,g8095,g7942,g2164,g6718,g2364,g2233,g9780,I16623,g10858,I13609,I10183,g6108,g11065,I7729,I5192,g2054,g6582,I14397,g8888,g7386,I11767,g4731,I8085,g2454,I5549,g8579,I12773,I13200,I10042,I12604,g7630,g8719,g4557,I9317,g2725,g2018,g1974,g8926,I11173,g4239,g4966,I8340,I14933,g7426,I14494,I11921,g11602,g8041,g8752,g8635,g6227,g5503,g4515,g7614,I12190,g10275,g4242,g10493,I16114,g4948,I7691,g9816,g1980,g4615,g11160,I13624,I17710,g6203,I9581,I15241,g4254,I16589,g10820,I16518,g8164,g7872,I15470,I5812,I17669,g2131,I7659,g3731,g7636,I6220,I4891,g8922,I8133,g8296,g2956,I15075,g8725,g8589,g3683,I6844,g11075,g2004,g10165,g10079,I17356,g8532,I13741,g7187,g2803,g4769,g5987,I11692,I11770,I17438,I9995,g5536,g6689,I17687,g10193,g10057,g10796,g5299,g4393,g5810,g10259,g7067,I6921,I15491,g8236,g10523,g11605,I7006,I13013,g8048,g5892,g6528,I17312,g2745,g2338,I5073,g8116,I11207,g6524,g7446,g3475,g3056,g11155,g3255,I15266,g7258,I12388,g7219,g8046,I14232,g7403,g3627,I6784,g4822,g3706,I12871,g6564,I16808,I11683,g11482,I8711,g2156,g2373,I12251,g7076,g10381,g2707,g2041,I8827,g4477,g10437,g10333,I5843,g4456,g4167,g7637,g10161,g3039,g2310,g3439,g7107,I12032,g6923,g8297,g10347,I8396,g4255,g3624,I11725,g5082,g4732,I11100,g5482,I14405,g8937,g10600,g4752,g8684,I13969,I8250,g5876,g2363,g6538,I13394,g10236,g4062,I7185,g2098,I4938,I9129,g7416,g4620,g10351,I15864,g10339,g6589,I10549,g3524,I15749,g2210,g11306,g7047,I7300,g2883,g11313,I17104,I12360,g7183,g4778,g10063,I17387,g11438,g8707,g8671,g6165,g10128,g6861,g5214,g10137,g6048,g9772,g6895,g2539,I5652,I6347,g6448,I10374,g9531,I14678,I15305,g6711,g6055,g11223,g11053,g9890,g6163,g3404,I9836,I9150,g6179,g9505,g9052,g9721,g2268,I13645,g4298,g3764,g8575,g8776,g4485,I8842,g6196,g7880,g7595,I12123,I11947,I17368,g8604,g8479,g10208,I16239,I17730,g8498,g6827,g4309,g9331,g7272,g8197,g10542,g11064,g7612,I12186,g2086,g7244,g7040,g7586,g2728,g7930,g6418,I11082,g7982,I12790,g4520,g5222,I17228,g11300,I17704,g4219,I10129,I6031,g4061,g10718,I6601,g3727,g7629,I15665,I11632,g2070,g3906,g11622,I13744,g10346,I15804,g5899,g4958,I10027,g10122,I7143,g10464,g10034,I15238,g6181,I11804,I14249,I17419,g6482,g10292,I15698,I9475,g5445,I9930,g6700,g11227,g6088,I10299,g7213,I11447,g2331,I16577,I8089,g2406,I13332,g8206,g4270,I11135,g6679,g4057,I15406,g11636,I12318,g11074,g10901,I11094,g11239,g11219,g4225,g2087,I17636,g3945,g2801,g2117,g5089,g4886,g3738,g3062,I14786,g9266,I12867,g9760,I6294,g11608,g3709,I6870,I7269,g4324,g2748,g6562,g10164,g7077,g10133,I9248,g5471,g4370,g2755,I16956,I7076,g2226,g2578,I10090,g6723,I10716,g8059,I10030,g8771,g11518,g6101,I9762,g7649,g2459,g4377,g6035,g3517,I6702,g10575,g7851,g11501,g3876,g8131,g10327,I15771,g2173,g7106,g4287,g6198,g7964,I12562,g8105,g7992,g2169,g8973,g10283,g2369,g6834,I7414,g5773,g4399,g6921,g2407,I14961,g9769,g1962,g2868,I8147,g6041,g2647,I13812,g5148,g6441,I13463,g8156,I14642,g3110,g11577,g7279,g5836,g4510,I12427,g7134,g2793,g4291,I12655,I17365,g10174,I15514,I16500,I16664,g10795,g9103,g2015,g6368,I13633,g3773,g7057,g4344,I5142,I7593,g4142,g7989,I15284,g7611,I12547,g11083,g11276,g10390,I16484,g10770,g9732,g5218,g11284,g5822,g4819,g3877,g9271,I12226,g8007,I7264,g3252,g2203,I15554,I10620,I5497,g2846,g7570,I13421,I16200,g10494,I5960,g4081,g8773,g6856,I10924,I10733,g5401,g8535,I7450,g8582,I13825,g7670,I17261,g3462,g4951,I8320,I11472,I16220,g5895,g7938,I8126,g3662,g4314,g5062,I13788,g10326,g4417,g7909,g2689,I12103,I11829,g6740,g10484,I16805,g10904,g8664,I15247,I10412,g5821,g7143,g9533,g8939,I13828,g2028,g8772,g10252,g8721,I10499,g10621,g7606,I12168,g2247,I5258,g4336,g2067,g2564,g7687,g4768,g11576,I17610,g6093,I13682,I6911,g2163,g6500,g10183,g5192,g4943,g3352,g11200,g3705,g10500,g11388,g4065,g2794,g3637,g4228,g4322,g5941,I14379,g4934,g4243,I11671,g6485,I10308,g8777,g6244,I13956,I6439,g5304,g3254,g9775,g11640,g3814,g5708,g5520,g11319,I13785,g3038,g1982,g4496,I7889,I8303,g4784,g5252,g7607,g11487,g5812,g3009,g9110,g6183,g2571,g5176,g6220,I5716,I5149,g10047,g4337,g4913,g11380,g2055,g10311,g2455,g9739,I6952,g9269,I9402,g5107,g7054,g4380,g1975,g7236,I11581,g2774,g3967,g3247,g11314,g7729,g5276,I15272,g9150,I9886,g7615,I12193,g6361,g4266,g4159,g9668,g2396,g10592,I9287,I17225,g11298,g7202,g5270,g4367,g7374,g6819,I12916,g11345,I7288,g2509,I16407,g10696,g2987,g5073,g10350,g11539,g6146,g7545,g2662,g5124,I9594,g7380,g6103,g5317,I11794,g8711,g7591,g8472,g4726,g2994,g5469,g7853,g4354,I7639,g7420,g5177,g8346,g11241,g10453,g6243,I5279,g6514,g7559,g8817,g10691,I16360,g8810,g8196,g6944,g8803,I6277,g6072,g8538,g2381,g9313,g10387,g4783,I7375,g2847,I5973,g6157,I12202,g6983,g8509,g8366,g9453,g4112,g7905,g7450,g4312,g4473,g6577,g10929,I12496,g7724,g5195,g6116,g2421,g4001,g3200,g8040,g10928,I9731,g5255,g5898,g6434,I10352,g4676,g5900,g5790,I5821,g2101,I11926,g6900,g8042,g4129,g5797,I9399,g4329,g4761,g11515,g11490,I7339,g7927,g8230,g6681,I11701,g5291,g3392,g6546,g3485,g2562,g6697,g5144,g4592,g6914,I11024,g11446,g6210,I12150,g6596,g4221,g8381,g2817,g3941,g7440,g8574,I10445,g5770,I17374,I11360,g8889,g7648,g5701,g4953,g3520,g10711,I6395,g2743,I15114,g9719,I17158,g11312,I16613,g11435,I6876,g5287,I16859,g3812,g5886,g11107,g6351,g10261,I13360,g8126,I17353,g3405,g9778,g4387,g9894,g8723,g8585,g4716,g6479,g3765,g3120,g5814,g5849,g3911,I16632,g9782,I5695,I5111,g6060,I16273,g10559,g5219,g4747,I10736,g4398,I13451,g10248,g2772,g2508,g7240,g8751,g4241,I9352,g5594,g9270,g8819,g9256,g6656,g6995,g7618,g3980,g2411,I5494,g10786,I13776,g4524,g3757,g5887,I9510,g10356,I15832,g5122,I17519,g6190,g2074,g4319,g6906,g10717,I16540,g4759,g3206,g5189,g4258,g4867,g6156,g4717,g2919,I10087,g9919,g2080,I14087,g8770,g2480,g6392,g6621,g5096,I11076,g2713,g6704,g11610,g4386,g10932,g4582,g5845,g4975,I7513,g11645,g5395,g5891,g11106,g4426,g10897,g6250,I10009,g4614,g9527,I14668,I7671,I12550,I7378,g6432,g7908,g7454,g8264,g6053,g9765,g11604,g9764,I16920,I16760,g3291,g2161,g7245,g6453,g4280,I7182,g4939,I11540,g6877,g2510,I15795,g3344,I16121,g6568,I7216,I12942,g4544,g3207,g2439,I7916,I12493,g2000,g8713,g11486,g2126,I6071,I14967,g7581,g10799,I15507,g3088,g4306,g7965,g5481,g4790,I9221,g1964,g10357,g7264,g10620,g10148,g11421,g4461,g6439,g4756,I17713,g8688,g8507,g7133,g10343,g8642,I14918,g4427,g8044,I15473,g10087,g8254,I6150,g11541,g11549,g9771,I12838,g2023,g11344,g4514,g5874,g5783,I9377,g4003,I6409,g5112,g7379,I8647,g11232,g5267,g11607,g6573,g9892,I8039,g3506,g3407,g4763,g7878,g8760,g11434,g4391,g6193,g3408,g3108,g2451,g7225,g6778,g7882,I17155,g4307,g4536,g10228,I15604,g4359,I13102,g8608,g8220,g7231,g4576,g3943,g4904,I10144,I14525,g8806,g11292,I16604,g6822,g4416,g7624,I14352,I5792,g10310,g7997,g2753,g4315,g3661,I15861,g6561,I11644,g10378,I15858,g5624,I11707,g6084,g8327,g8952,g4874,g6039,g5068,g6912,g3096,I11103,g3496,g6898,g8146,I5020,g5421,g8103,g7994,g3395,g2434,g3913,g6583,g6702,g4880,g5866,g8696,I7029,I14309,g8813,g2347,I7429,g10802,I7956,g7901,g4272,g10730,g7560,g6924,I17749,g8240,g5747,g4420,g5308,g7600,I12580,g7574,I6085,g10548,g11310,g3142,g6527,g4328,g11294,g3815,I11211,g5852,g6764,g2970,g6026,I11088,g9556,g10369,g10317,g3097,g5286,I6898,g6970,g2317,g4554,I15389,I15127,g3370,g5818,g8697,g8024,g10323,g11191,g2775,g3783,g5893,g5106,g8945,g3112,g3267,g7983,g4804,g6525,g2060,g6617,g6019,g6789,g8210,g5083,g3585,g11573,I5710,g5614,g7541,I7173,g7500,I13335,I9433,g3828,g10697,I16370,I9065,g4760,g11447,g8601,g2479,g10860,g2840,I10189,g7024,g10502,g2190,g4260,g2390,g11579,g7737,g3703,g4463,g7672,I12293,g6709,g11639,g9814,g5030,g6826,I14555,g2303,g8739,I12242,g4279,g9773,g11061,g10498,g9009,g6082,I9727,g4318,g4872,g7626,g5200,g4457,I8877,g6829,I17185,g10271,g9958,g4549,g7211,g11162,g5191,g3747,g10342,g3398,g6214,g10145,I9783,g5637,g7044,g2912,I13735,g8704,g4321,g10198,g5223,I7487,g7660,g8363,g10330,g10393,I7766,g10722,g6236,g11071,g8887,g11484,g11286,g6002,g11606,g11217,g10454,g4519,I7920,g5251,g6590,I11942,I12372,g7961,g6757,g4552,g4606,g6216,g8941,g10856,g7414,g3386,g4892,g7946,g3975,g4586,g7903,g2683,g3426,g5880,g6930,g8250,g2778,g5250,g5272,g7036,g9085,g4525,g7436,g8626,g6049,g8943,g10861,g11059,g2475,g8779,g3544,g11540,I6815,g5629,g5484,g6089,g7916,g11203,g5542,I8967,g7022,g3306,g2998,g3304,g6557,I12523,g3790,g4482,g6705,g5190,g6180,I15377,g9431,g9812,g3756,g4587,I12475,g5274,g4275,g4311,g3427,g5213,g8774,g10545,g10444,g10325,g7437,g8260,g4284,g8526,g6099,g3391,g10401,g5490,I14485,g11427,g5166,g6831,g4591,g6068,g7137,g7917,g9473,g10532,g1965,g4507,g6967,g6545,g2764,g11547,g7257,g6909,g8384,g7442,g8702,g2503,g11392,g10353,g3416,g6506,g8883,g3522,g11572,g2224,g6728,g10724,g2320,g4556,g3070,g3874,g8004,g2789,g5619,g5167,g11103,g2250,g9900,g11095,g4973,g7389,g7888,g7465,g4969,g8224,g2892,g5686,g10308,g4123,g8120,g6788,g5598,g4824,g9694,g10495,g2945,g11190,g8789,g8639,g9852,g9728,g9563,g5625,g4875,g9701,g7138,g10752,g11211,g11058,g11024,g8547,g8307,g10669,g7707,g4884,g3813,g4839,g9870,g6640,g9650,g9240,g5687,g7957,g3512,g7449,g4235,g4343,g11296,g9594,g9292,g9943,g9923,g9367,g5525,g8876,g10705,g10564,g9934,g9913,g9624,g6225,g6324,g10686,g6540,g8663,g11581,g6206,g3989,g7730,g7260,g7504,g7185,I5689,I5690,g7881,g11070,g9859,g9736,g9573,g8877,g11590,g2274,g6199,g8932,g5545,g5180,g5591,g8556,g8412,g11094,g5853,g5044,g6245,g4360,g8930,g5507,g11150,g3087,g8464,g8302,g9692,g4996,g7131,g11019,g9960,g9951,g9536,g11196,g11018,g10595,g10550,g10433,g10623,g10544,g4878,g5204,g4838,g8844,g8609,g6701,g6185,g10725,g5100,g4882,g8731,g5128,g6886,g8557,g8415,g8966,g8071,g11597,g9828,g9722,g9785,g2918,g9830,g9725,g8955,g9592,g5123,g7059,g6078,g7459,g11102,g7718,g7535,g9703,g5528,g5151,g9932,g9911,g5530,g2760,g8629,g6887,g6187,g6228,g5605,g6322,I6337,I6338,g8967,g5010,g3275,g2895,g7721,g9866,g9716,g10808,g10744,g3047,g4492,g3685,g8822,g8614,g10560,g11456,g9848,g9724,g9557,g4714,g6550,g5172,g10642,g3284,g2531,g9855,g5618,g6891,g7940,g11085,g4968,g8837,g8646,g9644,g9125,g5804,g8462,g8300,I6330,g11156,g6342,g9867,g9717,g4871,g10435,g7741,g9386,g9151,g8842,g8607,g9599,g9274,g8974,g5518,g9614,g9111,g4122,g7217,g4610,g11557,g2911,g11210,g7466,g9939,g9918,g11279,g10518,g10513,g10440,I16145,g8708,g7055,g5264,g6329,g8176,g8005,g7510,g4099,g3281,g11601,g11187,g6746,g6221,g8630,g9622,g11143,g10923,g9904,g9886,g9676,g8733,g6624,g11169,g8073,g9841,g9706,g9512,g5882,g5592,g8796,g8645,g11168,g4269,g5611,g8069,g9695,g10304,g8469,g8305,g4712,g6576,g5762,g10622,g11015,g5217,g5674,g9359,g9173,g9223,g8960,g11556,g9858,g5541,g4534,g5897,g6699,g6177,g6855,g3804,g3098,g5680,g9642,g5744,g8399,g9447,g9030,g11178,g8510,g8414,g6319,g11186,g3908,g2951,g6352,g9595,g9205,g4831,g4109,g5492,g8934,g10312,g6186,g9612,g9417,g9935,g9914,g8701,g10745,g10658,g11216,g9328,g8971,g11587,g6325,g7368,g6083,g6544,g5476,g7743,g4869,g5722,g6790,g5813,g8408,g10761,g7734,g8136,g7926,g5569,g9902,g9392,g8623,g5500,g2496,g6756,g3010,g5877,g8972,g6622,g11612,g9366,g11230,g4364,g9649,g5795,g5737,g4054,g6345,g5823,g11275,g9851,g6763,g5802,I16142,g10511,g10509,g10507,g9698,g4725,g9964,g9954,g5523,g8550,g8402,g8845,g8611,g2081,g6359,g11586,g11007,g5147,g5104,g5099,g4821,g5919,g5499,g4389,g3529,g6416,g3497,g4990,g9619,g9010,I6630,g6047,g9652,g10505,g10469,g9843,g9711,g9519,g5273,g11465,g4348,g11237,g9834,g9731,g6654,g5444,g3714,g11285,g9598,g8097,g8726,g6880,g4816,g3287,g10759,g9938,g9917,g10758,g10652,g9909,g9891,g7127,g6663,g11165,g6328,g8401,g11006,g5125,g4865,g4715,g4604,g2325,g5513,g11222,g6554,g7732,g9586,g5178,g4401,g4104,g4584,g7472,g11253,g9860,g8703,g11600,g9645,g11236,g4162,g3106,g6090,g9691,g11316,g11175,g8068,g9607,g9962,g9952,g6348,g9659,g9358,I6316,I6317,g4486,g9587,g8995,g5632,g8965,g4881,g11209,g8848,g8715,g4070,g3263,g6463,g8699,g7820,g11021,g5917,g6619,g6318,g6872,g11201,g10514,g10489,g4006,g9853,g11274,g8119,g9420,g5233,g7092,g6549,g11464,g4487,g2939,g7060,g6739,g5725,g11615,g2544,g11252,g5532,g11153,g3771,g9905,g9872,g9680,g7739,g6321,g8386,g8975,g2306,g6625,g7937,g8303,g8170,g5706,g2756,g8821,g8643,g10946,g5225,g4169,g5029,g11164,g4007,g4059,g4868,g5675,g4718,g10682,g6687,g7704,g4261,g3422,g5745,g8387,g7954,g11283,g8461,g8298,g10760,g11480,g6626,g8756,g6341,g10506,g9648,g7453,g5995,g6645,g5707,g7548,g11091,g11174,g8403,g8841,g8605,g6879,g8763,g4502,g9839,g9702,g9742,g6358,g5841,g5575,g8107,g10240,g11192,g9618,g5539,g8416,g9693,g11553,g7557,g5268,g9107,g10633,g7894,g8654,g9621,g6794,g5819,g4883,g3412,g7661,g2800,g3389,g3268,g9908,g3429,g6628,g5470,g7526,g2204,g5025,g6204,g4921,g4048,g8935,g2525,g9593,g4827,g10701,g10777,g10733,g8130,g9965,g9955,g3684,g11213,g5006,g9933,g9912,g8554,g8407,g9641,g6323,g10766,g10646,g6666,g4994,g5103,g11592,g3717,g6875,g9658,g6530,g6207,g8199,g7265,g9835,g9735,g6655,g3875,g7970,g7384,g5491,g8949,g11152,g9611,g6410,g2804,g10451,g4397,g7224,g5398,g5602,g6884,g8698,g8964,g11413,g4950,g5535,g7277,g6772,g8463,g8301,g2511,g10728,g6618,g6235,g6355,g4723,g3626,g8720,g6693,g11020,g11583,g8118,g8167,g7892,g8652,g5721,g10367,g10362,g9901,g6792,g11282,g7945,g11302,g11105,g3634,g8598,g8471,g7140,g9600,g9864,g11613,g5188,g7435,g7876,g4058,g6776,g5809,g10301,g4505,g9623,g10739,g11027,g10738,g8687,g8558,g6360,g9871,g5108,g11248,g4992,g11552,g9651,g11204,g7824,g5115,g8710,g7102,g9384,g2561,g9838,g9700,g9754,g3718,g10661,g10594,g11321,g8879,g7621,g8962,g10715,g2272,g8659,g9643,g8957,g5538,g4000,g4126,g4400,g4088,I5886,I5887,g6238,g10727,g8174,g5067,g5418,g10297,g6353,g11026,g11212,g6744,g4828,g10671,g4383,g2517,g5256,g4297,g4220,g8380,g8252,g7071,g9613,g8933,g5181,g7948,g11149,g9862,g11387,g7955,g4161,g11148,g2321,g9712,g8931,g11097,g3819,g11104,g2963,g6092,g4999,g7409,g4976,g6858,g4103,I6309,g6580,g5944,g5631,g9414,g9660,g9946,g9926,I6331,g9903,g9885,g9673,g10625,g6623,g11228,g11011,g6889,g7523,g7822,g8123,g11582,g4316,g3400,g10969,g3625,g5041,g9335,g9831,g9727,g9422,g8648,g4588,g8511,g8875,g5168,g7895,g7503,g8655,g3396,g4914,g9947,g9927,g5772,g5531,g5036,g10503,g8010,g7738,g8410,g6231,g5608,g10581,g10450,g10364,g2132,g2379,g4820,g9653,g10818,g8172,g10429,g5074,g9869,g10741,g10635,g8693,g5480,g4581,g3766,g2981,g8555,g8409,g9364,g8994,g11299,g6592,g7958,g4995,g4079,g2264,g2160,g3257,I6310,g5000,g3301,I5084,g9412,g9389,g10706,g10567,g10366,g10447,g10446,g10533,g5220,g10624,g10300,g5023,g4432,g4053,g7596,g5588,g6074,g9963,g9953,g3772,g3089,g5051,g8724,g4157,g9707,g8878,g10763,g10639,g6777,g8109,g7898,g7511,g11271,g11461,g5732,g11145,g11031,g9865,g9715,g9604,g8799,g8647,g11198,g6873,g6632,g6095,g9833,g9729,g6102,g7819,g11280,g7088,g9584,g9896,g8209,g6752,g11161,g8947,g5681,g7951,g9419,g5533,g8936,g10670,g11087,g4949,g6364,g5851,g7825,g10667,g7136,g6532,g9385,g9897,g9425,g3383,g5601,g7943,g11171,I6631,g7230,g6064,g4952,g8736,g6787,g8968,g10306,g11459,g11458,g5739,g7496,g4986,g11010,g5187,g3999,g8175,g8722,g5590,g7891,g7471,g8651,g5479,g11599,g6684,g6745,g6639,g3696,g4503,g6791,g8180,g4224,g5501,g8838,g8602,g10666,g11158,g9602,g5704,g4617,g3879,g9868,g11295,g11144,g9718,g3434,g4987,g6098,g9582,g3533,g8104,g9415,g8499,g8377,g9664,g2534,g8754,g9413,g6162,g3584,g4991,g6362,g5846,g10685,g11023,g7598,g11224,g11571,g4959,g5626,g9940,g9920,g4876,g6730,g9689,g10762,g6070,g9428,g9430,g8927,g7068,g8014,g7740,g11278,g5782,g9910,g4236,g11559,g9609,g11558,g6087,g4877,g10751,g10772,g10655,g8135,g11544,g5084,g8382,g10230,g7241,g3942,g10638,g4064,g9365,g9861,g9738,g9579,g8749,g11255,g11189,g10510,g2917,g11188,g9846,g7818,g11460,g11030,g11093,g7893,g7478,g8653,g10442,g6535,g8102,I5085,g3912,g7186,g4489,g9662,g9418,g11218,g10746,g10643,g7125,g7821,g6246,g8963,g7533,g10237,g7939,g8786,g8638,g10684,g11455,g8364,g2990,g9847,g7584,g5617,g5981,g5789,g4009,g11277,g6940,g6472,g7061,g6760,g11595,g5771,g8553,g8405,g4836,g5547,g4967,g6671,g7200,g7046,g4229,g8389,g6430,g8706,g4993,g6247,g11170,g7145,g5738,g3998,g6741,g11167,g11194,g11589,g4431,g7536,g9585,g2957,g11588,g5690,g6883,g4837,g8791,g8641,g6217,g11022,g5915,g4168,g8759,g5110,g11254,g7567,g4392,g3273,g9856,g9411,g5002,g11101,g11177,g11560,g8098,g3970,g4941,g6662,g7935,g6067,g9863,g9740,g6994,g6758,g4252,g11166,g7130,g11009,g5179,g7542,g11008,g5171,g3516,g7573,g3987,g11555,g9857,g9734,g9569,g8728,g8730,g8185,g8385,g7902,g4073,g8070,g5731,g11238,g8470,g8308,g5489,g3991,g7823,g4069,g11176,g11092,g11154,g9608,g11637,g2091,g8406,g5254,g8612,g9588,g8801,g8742,g7063,g10303,g5009,g9665,g8748,g11215,g10750,g5769,g3818,g8755,g6673,g7720,g4609,g7547,g7971,g11288,g7599,g6058,g6743,g4106,g6890,g7549,g7269,g8169,g11304,g9944,g9924,g7592,g8718,g8616,g9316,g7625,g8793,g8644,g2940,g11624,g10949,g2947,g4870,g3563,g10948,g2223,g8246,g7846,g5788,g4008,g9596,g5249,g11585,g4972,g11554,g7096,g10673,g4806,g2493,g9936,g9915,g2910,g9317,g10933,g10853,g8388,g8177,g7141,g10508,g4230,g10634,g9601,g9192,g6326,g7710,g8028,g7375,g5640,g5031,g4550,g7879,g7962,g9597,g5005,g6423,g8108,g5911,g3322,g9937,g9916,g9840,g9704,g9747,g10723,g8217,g11013,g5209,g9390,g11214,g6327,g5796,g5473,g6346,g5038,g6633,g11005,g5119,g8365,g7558,g4481,g4097,g7588,g4497,g9942,g9922,g6696,g10731,g5118,g10665,g8827,g8552,g5540,g4960,g8846,g8615,g5983,g6240,g7931,g11100,g11235,g5199,g6316,g7515,g5781,g8018,g7742,g2950,g5510,g6347,g9357,g11407,g10743,g5259,g5694,g10769,g11584,g4932,g10768,g10649,g4068,g6317,g5215,g4276,g4866,g6775,g10662,g8101,g5825,g3204,g5318,g7884,g7457,g3974,g9949,g9929,g10778,g7524,g6079,g7235,g9603,g9850,g9726,g9560,g7988,g5228,g5587,g5934,g8168,g9583,g10672,g8627,g8309,g10449,g10420,g11273,g8734,g5913,g4572,g6363,g11463,g8074,g8474,g8383,g11234,g4483,g11491,g5097,g5726,g5497,g7933,g9617,g9906,g9873,g9683,g11012,g5196,g7050,g10971,g10849,g8400,g4345,g9945,g9925,g7271,g5028,g9709,g4223,g10716,g10497,g11247,g6661,g11173,g6075,g8023,g7367,g9907,g9888,g9686,g10582,g5746,g9959,g9950,g7674,g9690,g5703,g4522,g4115,g7075,g10627,g4047,g2944,g6646,g7132,g11029,g7572,g8127,g7209,g11028,g10742,g8880,g10681,g9663,g5349,g8732,g3807,g8753,g5848,g3860,g8508,g8411,g8072,g5699,g11240,g6616,g6105,g10690,g7582,g9590,g4128,g6404,g6647,g10504,g9657,g4542,g5524,g9899,g7736,g10626,g6320,g7623,g10299,g7889,g10298,g8413,g3979,g5211,g4512,g7722,g9844,g9714,g9522,g4823,g5993,g5026,g8705,g10737,g10232,g6771,g5170,g8117,g9966,g9956,g5280,g7139,g11099,g6892,g9705,g10512,g11098,g8628,g5544,g11272,g5483,g9948,g9928,g4063,g11462,g6738,g7593,g11032,g10445,g8882,g10316,g5756,g4720,g9409,g8929,g6876,g4989,g9836,g9737,g6061,g8268,g6465,g5003,g9967,g9957,g5145,g4834,g4971,g10753,g5695,g7613,g10736,g11220,g7444,g4670,g4253,g8163,g7960,g10764,g5757,g10365,g8032,g7385,g11591,g2988,g7583,g11147,g5522,g9837,g9697,g9751,g9620,g11151,g11172,g7885,g5595,g5537,g9842,g9708,g9516,g4141,g4341,g7679,g7378,g5612,g3939,g7135,g10970,g11025,g9854,g9730,g9566,g7182,g9941,g9921,g6194,g4962,g4358,g8683,g4803,g8549,g5224,g8778,g11281,g8735,g11146,g3904,g2948,g8075,g9829,g9723,g7184,g11246,g6350,g5837,g5902,g2555,g6438,g5512,g5090,g7719,g3695,g7587,g9610,g3536,g8881,g4559,g10561,g10549,g5698,g11226,g10295,g5260,g10680,g11551,g11538,g9849,g5279,g8404,g5720,g8764,g11318,g11297,g9898,g9510,g7963,g9759,g9803,g6124,I14585,I5600,g9489,g3107,g2167,g9362,I14866,g4997,g10291,g9669,g6122,g9509,g5227,I15054,g5555,g10376,g8249,I15210,g9882,I5805,g2102,g2099,g2096,g2088,I15039,g8259,g10805,I15214,I15215,g8322,g9750,g8248,g8154,I6351,g2405,g2389,g2380,g2372,I16427,I14776,g4052,g2862,g2515,I14858,I15209,g2528,g2522,g9515,g3118,g2180,I5571,g2514,I5599,g9528,I5629,g2315,I5363,g8159,g10521,I16148,I16149,g8417,I14855,I15205,g9878,I15051,g9615,g8823,g8148,g2863,g2516,g9511,g9654,I15224,I15225,g8253,g9416,I15171,I15172,g9410,I15204,I14596,g9655,g10472,g10470,g10468,g10467,g10386,g10384,g10476,g10474,g8158,g9656,g9746,I5357,g9758,I5626,I15057,I15219,I15220,g9616,I14862,g2521,I14751,g9591,g9757,g9815,I14835,I16161,g10479,g10478,g10477,g10475,g2353,g9776,I5804,I15199,g8153,g9881,g9426,g9423,g8262,g2499,I5570,I14607,g9388,g10807,I16160,g10394,g10392,g10482,g10481,I15042,g9589,g9667,I14827,g9779,g9391,g2309,I5358,I15177,g9876,g9421,g5186,I6350,g8162,I14779,g2305,I5351,I5352,I15176,g9879,g10562,g9606,I14822,I15200,g9880,I14582,g8247,I5576,g4476,g2538,I5649,g9605,g9781,g9363,I14831,g8263,g9361,g5780,I15048,g9647,g9817,I14602,I15033,g2445,g2437,g2433,g2419,I5366,g9506,g8161,g2316,g4675,g9387,I15045,g9808,g2501,g9877,g10529,g9874,g8157,g6899,g9646,g2111,g2109,g2106,g2104,I5612,I5613,I5593,I5591,g8970,g8839,I10519,I11279,I11278,g3978,I5264,I5263,I8640,g4278,I6761,g2943,I6760,I17400,g11418,g11416,I5450,I5449,I16060,g10372,I16058,I6746,g2938,I11975,I11973,I12136,I11937,I11935,g2959,I6167,I6168,I5878,g2120,g2115,I5619,I5620,g5552,I6468,I6467,I8796,g4672,I8795,I15891,I15892,I5611,g8738,I6716,I6714,I7685,g3460,I7683,I12108,I12106,I6747,g2236,I5230,I5231,I12075,I12076,I15870,g10358,I16067,I16065,I7562,I13531,I13529,I8797,I17584,I11936,I15257,I15256,I13505,I13506,g8824,g8502,g8501,I6186,g11496,I17504,I17505,I16001,I15999,I6125,g2215,I6124,I11909,I11907,I12040,I12038,I13909,I13907,I6771,I6772,I11908,I16008,I16009,I13908,I7034,I7035,I8650,I9947,I9948,I16066,g10428,I6144,I6145,I11242,I11241,I15993,I15994,I6187,g6027,I5500,I11974,I12062,I12060,I8771,I8772,I5184,I13293,I6200,I6199,I13265,I5024,I5023,I7863,I13991,I13992,I13660,I13661,I6143,I13990,I11510,I11508,g5034,I5229,I12047,I12045,I10771,I10769,I16045,I16046,I12061,I5104,I13530,I6447,I4956,I4954,I8481,g3530,I8479,I8739,I8740,I6880,I6879,I15431,I15430,I12020,I12019,I16331,I16332,I16469,I16467,I5014,I5013,I13523,I13521,I16039,I16037,I16468,I12046,I16038,g10427,I8676,g4374,I12113,I8761,g4616,g10422,I15992,I5036,I5034,I14263,g8843,I13249,I13250,I5135,I5485,I5486,I7033,I15443,I15441,I6166,I8624,g4267,I16015,g10425,I8677,I8576,g4234,I8575,I14613,g9204,I14612,I8716,g4601,I8715,I6715,I13514,I13515,I12003,I12002,g2177,I5127,I5128,I8577,I17395,g11414,I17393,I11280,I5265,I6989,I6988,I13274,I13272,I10507,I5164,I14443,I14444,I9559,I9557,I5592,I13077,I13078,I8717,I5296,I5295,I8625,I8626,I4911,I4912,I16000,g10423,I5371,I5185,I5186,I5675,I8544,g4218,I8543,I10520,I10521,I5297,I13537,I13283,g4749,I11982,I11980,I8514,g4873,I8513,I13091,I13089,I6126,I15908,g10302,I15906,I8763,g8825,g8506,I16007,g10424,I5865,g2107,g2105,I5604,I5517,I5518,I6111,I6109,I4929,I4930,I13522,I10770,I5539,I5538,I17394,g11415,I13553,I13552,I8642,I17296,I17297,I14278,I14279,I4910,I6794,I6792,I5484,I15442,I10931,I10932,I8779,I8780,g2354,I15615,g10043,g10153,I17281,I5470,I5468,I11509,I5025,I14272,I14270,I6208,I6209,I17290,I17288,I7563,I7564,I5006,I5005,I12128,I12126,I5105,I6323,I6322,I12093,I12094,I6666,g2776,I6664,g3623,I6762,I5373,I8529,I8527,I5283,I5282,I7224,I7223,I5007,I5459,I17295,I5015,I14264,I14265,I16073,I16072,g3205,I8652,I9558,I5203,I5202,I6806,I6807,I6469,I12145,I12143,I12127,I13302,I13300,I5502,I9574,I6448,I6449,I8670,I8669,I15453,I15451,I7876,I7875,I14203,I14202,I15607,g10149,g10144,I5324,I5325,I8738,g10434,g5859,I8606,I8604,I12087,I12085,I13248,I4979,I4980,I12069,I12067,g8942,I12068,I17503,I7877,I5165,I6289,I6287,I6777,I8562,I8563,I15890,I13090,g8006,g11474,I17460,I17461,I13513,I4986,I4987,I5204,I13504,I6207,I12086,I8545,I8180,I8178,I8591,I8589,I10930,I17402,I13294,I13295,I12144,g8757,g2961,I14211,I14209,I8515,I5316,I5317,I9946,I8750,g4613,I5605,I14204,I16051,g10371,g10373,g10360,g6037,I13858,I13859,I15872,I8528,g4879,I13901,I13902,g8542,I6838,I6836,I17307,I17305,g4538,I15452,I13857,I13765,I8671,g10370,I16044,g10363,g5360,I5106,I8804,g4677,I8803,I16016,I16017,I17487,I17485,I4995,I12092,I8678,I5126,I5372,I17306,I11995,I7225,I11261,g8545,I6110,I4942,I4941,I15899,I15900,g5527,g10443,g5350,I16081,g10374,I16079,I8641,I6178,I6176,I12074,I5451,I7322,I7323,I6288,I8179,I6805,I17486,I4928,g10286,I16330,I9575,I13887,I13886,I8787,I8788,I5315,g10285,I13869,I13867,I13868,I13259,I13258,g3261,I16074,I5136,I5137,I5460,I5461,I8605,I6770,g11449,I17401,g11448,I15717,g10231,I15716,I14210,I17569,I17567,I13878,I13876,I5606,I14442,I11996,I11997,I14277,I17568,I7321,I6990,g8847,I9006,I4985,I8651,I13545,I13544,I13894,I13895,I6138,I6136,I13076,g2205,I13260,I5501,I17586,I13900,I6201,I14217,g8826,I14216,I9007,I13561,I13559,g10229,I17493,I17492,I12215,I12214,I11262,I11263,I6225,I6226,I13309,I13307,I5676,I5677,I6826,I6827,I13308,g8190,g2792,I5879,I5880,g3061,I17585,I6881,I12138,I8729,g4605,I8728,I15871,I5866,I5867,I6793,I6487,I16080,I13893,I12115,I6748,I6224,I8805,I15880,I15878,I16031,I16030,I14271,I13267,I15616,I15617,I4966,I4964,I8752,I15432,g10438,g6032,g3011,I8480,I16087,I16086,g3734,I14218,I4955,I8786,g4639,g10480,I11915,I11914,I8770,g4619,I5516,g8541,I6188,I5892,I5891,I13766,I13767,I15258,I13266,I6825,I17283,g5277,I5035,g10375,I15879,g10359,I12114,I12107,g2500,g10430,g5999,I13285,I13877,g2795,I5893,I13560,g4259,I5166,I14614,I4965,I4943,I16023,g10426,I16059,g8737,I9576,I16052,I16053,I12004,g5573,I6837,I8730,I4978,I6177,I17051,I7864,I7865,I6665,I12216,I13554,g10368,I13284,I6137,I5529,I5530,I17282,I5618,I8664,I8662,I11916,g7717,I4972,I4971,I13273,I10509,I10508,I6778,I6779,I5469,g4251,I13546,I4996,I4997,I13539,I16032,I5323,I13538,I5540,I8778,g4286,I17052,I17053,g10287,I15898,g7978,g4227,I8561,I8762,I8751,I15907,I4973,I16024,I16025,g4455,I5342,I5341,I12137,g10483,I16088,I17289,g4630,I15609,I15608,g10436,g6023,I17459,I13301,I11981,I8663,I15718,I5284,g4607,g8840,g10441,g5345,g10432,g5938,I12021,I6489,I5528,I13659,I5343,I12039,I9008,I6488,I13888,I17494,I7684,g3221,I6324,I8590,I11243,g10324,g10239,g4974,g10322;
AND2X1 AND1 (.Y(CK2), .A(CK), .B(CK));
INVX1 INV1 (.Y(SE_B), .A(SE));
AND2X1 AND2 (.Y(CK1), .A(CK), .B(SE_B));
DFFX1 DFF_17 (.CK(CK1), .D(g7354), .Q(g1574));
DFFX1 DFF_18 (.CK(CK1), .D(g7816), .Q(g1864));
DFFX1 DFF_19 (.CK(CK1), .D(g11439), .Q(g369));
DFFX1 DFF_20 (.CK(CK1), .D(g7356), .Q(g1580));
NAND2X1 AND2_690 (.Y(g5257),.A(g691),.B(g4755));
NAND2X1 AND2_691 (.Y(g4732),.A(g391),.B(g3372));
AND2X1 AND2_692 (.Y(g3108),.A(I6330),.B(I6331));
AND2X1 AND2_696 (.Y(g5605),.A(g4828),.B(g704));
NAND2X1 AND2_697 (.Y(g6623),.A(g55),.B(g6170));
AND2X1 AND2_698 (.Y(g11228),.A(g466),.B(g11060));
AND2X1 AND2_699 (.Y(g11011),.A(g1968),.B(g10809));
NAND2X1 AND2_700 (.Y(g6889),.A(g1941),.B(g6427));
AND2X1 AND2_701 (.Y(g8040),.A(g7523),.B(g5128));
DFFX1 DFF_21 (.CK(CK1), .D(g6846), .Q(g1736));
DFFX1 DFF_22 (.CK(CK1), .D(g10774), .Q(g39));
DFFX1 DFF_23 (.CK(CK1), .D(g11182), .Q(g1651));
DFFX1 DFF_24 (.CK(CK1), .D(g7330), .Q(g1424));
DFFX1 DFF_25 (.CK(CK1), .D(g1736), .Q(g1737));
DFFX1 DFF_26 (.CK(CK1), .D(g11037), .Q(g1672));
DFFX1 DFF_27 (.CK(CK1), .D(g6805), .Q(g1077));
DFFX1 DFF_28 (.CK(CK1), .D(g8279), .Q(g1231));
INVX1 NOT_4936 (.Y(I16114),.A(g10387));
INVX1 NOT_4937 (.Y(g4783),.A(g3829));
INVX1 NOT_4938 (.Y(g6043),.A(I9662));
INVX1 NOT_4939 (.Y(I12910),.A(g7922));
INVX1 NOT_4940 (.Y(I7375),.A(g4062));
INVX1 NOT_4941 (.Y(g2847),.A(I5973));
INVX1 NOT_4942 (.Y(g8780),.A(I14077));
INVX1 NOT_4943 (.Y(g6443),.A(g6157));
INVX1 NOT_4944 (.Y(I12202),.A(g6983));
INVX1 NOT_4945 (.Y(g8509),.A(g8366));
INVX1 NOT_4946 (.Y(g9453),.A(g9100));
INVX1 NOT_4947 (.Y(g4112),.A(g2994));
INVX1 NOT_4948 (.Y(g7905),.A(g7450));
DFFX1 DFF_29 (.CK(CK1), .D(g8079), .Q(g4));
DFFX1 DFF_30 (.CK(CK1), .D(g7785), .Q(g774));
DFFX1 DFF_31 (.CK(CK1), .D(g6815), .Q(g1104));
DFFX1 DFF_32 (.CK(CK1), .D(g7290), .Q(g1304));
DFFX1 DFF_33 (.CK(CK1), .D(g7325), .Q(g243));
DFFX1 DFF_51 (.CK(CK1), .D(g11333), .Q(g496));
DFFX1 DFF_52 (.CK(CK1), .D(g11472), .Q(g981));
DFFX1 DFF_53 (.CK(CK1), .D(g4896), .Q(g878));
DFFX1 DFF_54 (.CK(CK1), .D(g5653), .Q(g590));
DFFX1 DFF_55 (.CK(CK1), .D(g4182), .Q(g829));
DFFX1 DFF_56 (.CK(CK1), .D(g6811), .Q(g1095));
DFFX1 DFF_57 (.CK(CK1), .D(g9344), .Q(g704));
DFFX1 DFF_58 (.CK(CK1), .D(g7302), .Q(g1265));
DFFX1 DFF_59 (.CK(CK1), .D(g7814), .Q(g1786));
AND2X1 AND2_693 (.Y(g4753),.A(g481),.B(g3386));
AND2X1 AND2_694 (.Y(g9903),.A(g9885),.B(g9673));
AND2X1 AND2_695 (.Y(g10625),.A(g10546),.B(g4552));
DFFX1 DFF_60 (.CK(CK1), .D(g8429), .Q(g682));
DFFX1 DFF_61 (.CK(CK1), .D(g7292), .Q(g1296));
DFFX1 DFF_62 (.CK(CK1), .D(g6295), .Q(g587));
DFFX1 DFF_63 (.CK(CK1), .D(g7777), .Q(g52));
DFFX1 DFF_64 (.CK(CK1), .D(g8065), .Q(g646));
DFFX1 DFF_65 (.CK(CK1), .D(g5649), .Q(g327));
DFFX1 DFF_66 (.CK(CK1), .D(g6836), .Q(g1389));
DFFX1 DFF_67 (.CK(CK1), .D(g7311), .Q(g1371));
DFFX1 DFF_68 (.CK(CK1), .D(g1955), .Q(g1956));
DFFX1 DFF_69 (.CK(CK1), .D(g11038), .Q(g1675));
DFFX1 DFF_70 (.CK(CK1), .D(g11508), .Q(g354));
DFFX1 DFF_71 (.CK(CK1), .D(g7285), .Q(g113));
DFFX1 DFF_72 (.CK(CK1), .D(g8063), .Q(g639));
DFFX1 DFF_73 (.CK(CK1), .D(g11041), .Q(g1684));
DFFX1 DFF_74 (.CK(CK1), .D(g8448), .Q(g1639));
DFFX1 DFF_75 (.CK(CK1), .D(g8080), .Q(g1791));
DFFX1 DFF_76 (.CK(CK1), .D(g7323), .Q(g248));
DFFX1 DFF_77 (.CK(CK1), .D(g4907), .Q(g1707));
DFFX1 DFF_78 (.CK(CK1), .D(g5668), .Q(g1759));
DFFX1 DFF_79 (.CK(CK1), .D(g11507), .Q(g351));
DFFX1 DFF_80 (.CK(CK1), .D(g1956), .Q(g1957));
DFFX1 DFF_81 (.CK(CK1), .D(g7364), .Q(g1604));
DFFX1 DFF_93 (.CK(CK1), .D(g878), .Q(g876));
DFFX1 DFF_94 (.CK(CK1), .D(g6808), .Q(g1086));
DFFX1 DFF_95 (.CK(CK1), .D(g8444), .Q(g1486));
DFFX1 DFF_96 (.CK(CK1), .D(g10881), .Q(g1730));
DFFX1 DFF_97 (.CK(CK1), .D(g7328), .Q(g1504));
DFFX1 DFF_98 (.CK(CK1), .D(g8440), .Q(g1470));
DFFX1 DFF_99 (.CK(CK1), .D(g8437), .Q(g822));
DFFX1 DFF_100 (.CK(CK1), .D(g6291), .Q(g583));
DFFX1 DFF_101 (.CK(CK1), .D(g11039), .Q(g1678));
DFFX1 DFF_102 (.CK(CK1), .D(g8423), .Q(g174));
DFFX1 DFF_103 (.CK(CK1), .D(g7810), .Q(g1766));
DFFX1 DFF_104 (.CK(CK1), .D(g8450), .Q(g1801));
DFFX1 DFF_105 (.CK(CK1), .D(g7317), .Q(g186));
DFFX1 DFF_106 (.CK(CK1), .D(g11403), .Q(g959));
DFFX1 DFF_107 (.CK(CK1), .D(g6314), .Q(g1169));
DFFX1 DFF_108 (.CK(CK1), .D(g7806), .Q(g1007));
DFFX1 DFF_109 (.CK(CK1), .D(g8993), .Q(g1407));
DFFX1 DFF_110 (.CK(CK1), .D(g7794), .Q(g1059));
DFFX1 DFF_111 (.CK(CK1), .D(g7817), .Q(g1868));
DFFX1 DFF_112 (.CK(CK1), .D(g6797), .Q(g758));
DFFX1 DFF_113 (.CK(CK1), .D(g6337), .Q(g1718));
DFFX1 DFF_114 (.CK(CK1), .D(g11265), .Q(g396));
DFFX1 DFF_115 (.CK(CK1), .D(g7808), .Q(g1015));
DFFX1 DFF_116 (.CK(CK1), .D(g10872), .Q(g38));
DFFX1 DFF_117 (.CK(CK1), .D(g5655), .Q(g632));
DFFX1 DFF_118 (.CK(CK1), .D(g7335), .Q(g1415));
DFFX1 DFF_119 (.CK(CK1), .D(g8278), .Q(g1227));
DFFX1 DFF_120 (.CK(CK1), .D(g10878), .Q(g1721));
DFFX1 DFF_121 (.CK(CK1), .D(g883), .Q(g882));
DFFX1 DFF_122 (.CK(CK1), .D(g4906), .Q(g16));
DFFX1 DFF_123 (.CK(CK1), .D(g7767), .Q(g284));
DFFX1 DFF_124 (.CK(CK1), .D(g11256), .Q(g426));
DFFX1 DFF_125 (.CK(CK1), .D(g7310), .Q(g219));
DFFX1 DFF_126 (.CK(CK1), .D(g1360), .Q(g1216));
DFFX1 DFF_127 (.CK(CK1), .D(g7289), .Q(g806));
DFFX1 DFF_128 (.CK(CK1), .D(g8992), .Q(g1428));
DFFX1 DFF_129 (.CK(CK1), .D(g6287), .Q(g579));
DFFX1 DFF_130 (.CK(CK1), .D(g7351), .Q(g1564));
DFFX1 DFF_131 (.CK(CK1), .D(g5662), .Q(g1741));
DFFX1 DFF_132 (.CK(CK1), .D(g7309), .Q(g225));
DFFX1 DFF_133 (.CK(CK1), .D(g7766), .Q(g281));
DFFX1 DFF_134 (.CK(CK1), .D(g11627), .Q(g1308));
DFFX1 DFF_135 (.CK(CK1), .D(g9930), .Q(g611));
DFFX1 DFF_136 (.CK(CK1), .D(g5654), .Q(g631));
DFFX1 DFF_137 (.CK(CK1), .D(g9823), .Q(g1217));
DFFX1 DFF_138 (.CK(CK1), .D(g7359), .Q(g1589));
DFFX1 DFF_139 (.CK(CK1), .D(g8439), .Q(g1466));
DFFX1 DFF_140 (.CK(CK1), .D(g7353), .Q(g1571));
DFFX1 DFF_141 (.CK(CK1), .D(g7815), .Q(g1861));
DFFX1 DFF_142 (.CK(CK1), .D(g7307), .Q(g1365));
DFFX1 DFF_143 (.CK(CK1), .D(g11594), .Q(g1448));
DFFX1 DFF_144 (.CK(CK1), .D(g6335), .Q(g1711));
DFFX1 DFF_145 (.CK(CK1), .D(g6309), .Q(g1133));
DFFX1 DFF_146 (.CK(CK1), .D(g11635), .Q(g1333));
DFFX1 DFF_147 (.CK(CK1), .D(g8426), .Q(g153));
DFFX1 DFF_148 (.CK(CK1), .D(g11404), .Q(g962));
DFFX1 DFF_149 (.CK(CK1), .D(g6799), .Q(g766));
DFFX1 DFF_150 (.CK(CK1), .D(g6296), .Q(g588));
DFFX1 DFF_151 (.CK(CK1), .D(g11331), .Q(g486));
DFFX1 DFF_152 (.CK(CK1), .D(g11469), .Q(g471));
DFFX1 DFF_153 (.CK(CK1), .D(g7322), .Q(g1397));
DFFX1 DFF_154 (.CK(CK1), .D(g6288), .Q(g580));
DFFX1 DFF_155 (.CK(CK1), .D(g8288), .Q(g1950));
DFFX1 DFF_156 (.CK(CK1), .D(g755), .Q(g756));
DFFX1 DFF_157 (.CK(CK1), .D(g5656), .Q(g635));
DFFX1 DFF_158 (.CK(CK1), .D(g6814), .Q(g1101));
DFFX1 DFF_159 (.CK(CK1), .D(g11044), .Q(g549));
DFFX1 DFF_160 (.CK(CK1), .D(g7788), .Q(g1041));
DFFX1 DFF_161 (.CK(CK1), .D(g11180), .Q(g105));
DFFX1 DFF_162 (.CK(CK1), .D(g11036), .Q(g1669));
DFFX1 DFF_163 (.CK(CK1), .D(g7308), .Q(g1368));
DFFX1 DFF_164 (.CK(CK1), .D(g7340), .Q(g1531));
DFFX1 DFF_165 (.CK(CK1), .D(g7327), .Q(g1458));
DFFX1 DFF_166 (.CK(CK1), .D(g10877), .Q(g572));
DFFX1 DFF_167 (.CK(CK1), .D(g7805), .Q(g1011));
DFFX1 DFF_168 (.CK(CK1), .D(g10867), .Q(g33));
DFFX1 DFF_169 (.CK(CK1), .D(g7331), .Q(g1411));
DFFX1 DFF_170 (.CK(CK1), .D(g6813), .Q(g1074));
DFFX1 DFF_171 (.CK(CK1), .D(g11259), .Q(g444));
DFFX1 DFF_172 (.CK(CK1), .D(g8441), .Q(g1474));
DFFX1 DFF_173 (.CK(CK1), .D(g6806), .Q(g1080));
DFFX1 DFF_174 (.CK(CK1), .D(g6336), .Q(g1713));
DFFX1 DFF_175 (.CK(CK1), .D(g5651), .Q(g333));
DFFX1 DFF_176 (.CK(CK1), .D(g7762), .Q(g269));
DFFX1 DFF_177 (.CK(CK1), .D(g11266), .Q(g401));
DFFX1 DFF_178 (.CK(CK1), .D(g11409), .Q(g1857));
DFFX1 DFF_179 (.CK(CK1), .D(g7336), .Q(g9));
DFFX1 DFF_180 (.CK(CK1), .D(g8782), .Q(g664));
DFFX1 DFF_181 (.CK(CK1), .D(g11405), .Q(g965));
DFFX1 DFF_182 (.CK(CK1), .D(g7324), .Q(g1400));
DFFX1 DFF_183 (.CK(CK1), .D(g5652), .Q(g309));
DFFX1 DFF_184 (.CK(CK1), .D(g8077), .Q(g814));
DFFX1 DFF_185 (.CK(CK1), .D(g7319), .Q(g231));
DFFX1 DFF_186 (.CK(CK1), .D(g11048), .Q(g557));
DFFX1 DFF_187 (.CK(CK1), .D(g6294), .Q(g586));
DFFX1 DFF_188 (.CK(CK1), .D(g875), .Q(g869));
DFFX1 DFF_189 (.CK(CK1), .D(g7316), .Q(g1383));
DFFX1 DFF_190 (.CK(CK1), .D(g8425), .Q(g158));
DFFX1 DFF_191 (.CK(CK1), .D(g5657), .Q(g627));
DFFX1 DFF_192 (.CK(CK1), .D(g7799), .Q(g1023));
DFFX1 DFF_193 (.CK(CK1), .D(g7755), .Q(g259));
DFFX1 DFF_194 (.CK(CK1), .D(g1206), .Q(g1361));
DFFX1 DFF_195 (.CK(CK1), .D(g11633), .Q(g1327));
DFFX1 DFF_196 (.CK(CK1), .D(g8067), .Q(g654));
DFFX1 DFF_197 (.CK(CK1), .D(g7770), .Q(g293));
DFFX1 DFF_198 (.CK(CK1), .D(g11656), .Q(g1346));
DFFX1 DFF_199 (.CK(CK1), .D(g8873), .Q(g1633));
DFFX1 DFF_200 (.CK(CK1), .D(g5666), .Q(g1753));
DFFX1 DFF_201 (.CK(CK1), .D(g7329), .Q(g1508));
DFFX1 DFF_202 (.CK(CK1), .D(g7297), .Q(g1240));
DFFX1 DFF_203 (.CK(CK1), .D(g11326), .Q(g538));
DFFX1 DFF_204 (.CK(CK1), .D(g11269), .Q(g416));
DFFX1 DFF_205 (.CK(CK1), .D(g11325), .Q(g542));
DFFX1 DFF_206 (.CK(CK1), .D(g11040), .Q(g1681));
S_DFFX1 S_DFF_207 (.CK(CK2), .D(g11440), .SE(SE), .SI(SI), .Q(g374));
S_DFFX1 S_DFF_208 (.CK(CK2), .D(g11050), .SE(SE), .SI(g374), .Q(g563));
S_DFFX1 S_DFF_209 (.CK(CK2), .D(g8284), .SE(SE), .SI(g563), .Q(g1914));
S_DFFX1 S_DFF_210 (.CK(CK2), .D(g11328), .SE(SE), .SI(g1914), .Q(g530));
S_DFFX1 S_DFF_211 (.CK(CK2), .D(g11052), .SE(SE), .SI(g530), .Q(g575));
S_DFFX1 S_DFF_212 (.CK(CK2), .D(g9355), .SE(SE), .SI(g575), .Q(g1936));
S_DFFX1 S_DFF_213 (.CK(CK2), .D(g7778), .SE(SE), .SI(g1936), .Q(g55));
S_DFFX1 S_DFF_214 (.CK(CK2), .D(g6299), .SE(SE), .SI(g55), .Q(g1117));
S_DFFX1 S_DFF_215 (.CK(CK2), .D(g1356), .SE(SE), .SI(g1117), .Q(g1317));
S_DFFX1 S_DFF_216 (.CK(CK2), .D(g11509), .SE(SE), .SI(g1317), .Q(g357));
S_DFFX1 S_DFF_217 (.CK(CK2), .D(g11263), .SE(SE), .SI(g357), .Q(g386));
S_DFFX1 S_DFF_218 (.CK(CK2), .D(g7363), .SE(SE), .SI(g386), .Q(g1601));
S_DFFX1 S_DFF_219 (.CK(CK2), .D(g11046), .SE(SE), .SI(g1601), .Q(g553));
S_DFFX1 S_DFF_220 (.CK(CK2), .D(g7747), .SE(SE), .SI(g553), .Q(g166));
S_DFFX1 S_DFF_221 (.CK(CK2), .D(g11334), .SE(SE), .SI(g166), .Q(g501));
S_DFFX1 S_DFF_222 (.CK(CK2), .D(g7758), .SE(SE), .SI(g501), .Q(g262));
S_DFFX1 S_DFF_223 (.CK(CK2), .D(g8694), .SE(SE), .SI(g262), .Q(g1840));
S_DFFX1 S_DFF_224 (.CK(CK2), .D(g7783), .SE(SE), .SI(g1840), .Q(g70));
S_DFFX1 S_DFF_225 (.CK(CK2), .D(g5646), .SE(SE), .SI(g70), .Q(g318));
S_DFFX1 S_DFF_226 (.CK(CK2), .D(g6818), .SE(SE), .SI(g318), .Q(g1356));
S_DFFX1 S_DFF_227 (.CK(CK2), .D(g6800), .SE(SE), .SI(g1356), .Q(g794));
S_DFFX1 S_DFF_228 (.CK(CK2), .D(g10870), .SE(SE), .SI(g794), .Q(g36));
S_DFFX1 S_DFF_229 (.CK(CK2), .D(g7773), .SE(SE), .SI(g36), .Q(g302));
S_DFFX1 S_DFF_230 (.CK(CK2), .D(g11513), .SE(SE), .SI(g302), .Q(g342));
S_DFFX1 S_DFF_231 (.CK(CK2), .D(g7299), .SE(SE), .SI(g342), .Q(g1250));
S_DFFX1 S_DFF_232 (.CK(CK2), .D(g6301), .SE(SE), .SI(g1250), .Q(g1163));
S_DFFX1 S_DFF_233 (.CK(CK2), .D(g2044), .SE(SE), .SI(g1163), .Q(g1810));
S_DFFX1 S_DFF_234 (.CK(CK2), .D(g7800), .SE(SE), .SI(g1810), .Q(g1032));
S_DFFX1 S_DFF_235 (.CK(CK2), .D(g8990), .SE(SE), .SI(g1032), .Q(g1432));
S_DFFX1 S_DFF_236 (.CK(CK2), .D(g7792), .SE(SE), .SI(g1432), .Q(g1053));
S_DFFX1 S_DFF_237 (.CK(CK2), .D(g7326), .SE(SE), .SI(g1053), .Q(g1453));
S_DFFX1 S_DFF_238 (.CK(CK2), .D(g11511), .SE(SE), .SI(g1453), .Q(g363));
S_DFFX1 S_DFF_239 (.CK(CK2), .D(g5650), .SE(SE), .SI(g363), .Q(g330));
S_DFFX1 S_DFF_240 (.CK(CK2), .D(g6303), .SE(SE), .SI(g330), .Q(g1157));
S_DFFX1 S_DFF_241 (.CK(CK2), .D(g6330), .SE(SE), .SI(g1157), .Q(g1357));
S_DFFX1 S_DFF_242 (.CK(CK2), .D(g10869), .SE(SE), .SI(g1357), .Q(g35));
S_DFFX1 S_DFF_243 (.CK(CK2), .D(g8569), .SE(SE), .SI(g35), .Q(g928));
S_DFFX1 S_DFF_244 (.CK(CK2), .D(g7757), .SE(SE), .SI(g928), .Q(g261));
S_DFFX1 S_DFF_245 (.CK(CK2), .D(g11337), .SE(SE), .SI(g261), .Q(g516));
S_DFFX1 S_DFF_246 (.CK(CK2), .D(g7759), .SE(SE), .SI(g516), .Q(g254));
S_DFFX1 S_DFF_247 (.CK(CK2), .D(g8076), .SE(SE), .SI(g254), .Q(g778));
S_DFFX1 S_DFF_248 (.CK(CK2), .D(g4190), .SE(SE), .SI(g778), .Q(g861));
S_DFFX1 S_DFF_249 (.CK(CK2), .D(g8871), .SE(SE), .SI(g861), .Q(g1627));
S_DFFX1 S_DFF_250 (.CK(CK2), .D(g7293), .SE(SE), .SI(g1627), .Q(g1292));
S_DFFX1 S_DFF_251 (.CK(CK2), .D(g7769), .SE(SE), .SI(g1292), .Q(g290));
S_DFFX1 S_DFF_252 (.CK(CK2), .D(g5671), .SE(SE), .SI(g290), .Q(g1850));
S_DFFX1 S_DFF_253 (.CK(CK2), .D(g7288), .SE(SE), .SI(g1850), .Q(g770));
S_DFFX1 S_DFF_254 (.CK(CK2), .D(g7357), .SE(SE), .SI(g770), .Q(g1583));
S_DFFX1 S_DFF_255 (.CK(CK2), .D(g11468), .SE(SE), .SI(g1583), .Q(g466));
S_DFFX1 S_DFF_256 (.CK(CK2), .D(g7350), .SE(SE), .SI(g466), .Q(g1561));
S_DFFX1 S_DFF_257 (.CK(CK2), .D(g4899), .SE(SE), .SI(g1561), .Q(g1527));
S_DFFX1 S_DFF_258 (.CK(CK2), .D(g7345), .SE(SE), .SI(g1527), .Q(g1546));
S_DFFX1 S_DFF_259 (.CK(CK2), .D(g7768), .SE(SE), .SI(g1546), .Q(g287));
S_DFFX1 S_DFF_260 (.CK(CK2), .D(g11049), .SE(SE), .SI(g287), .Q(g560));
S_DFFX1 S_DFF_261 (.CK(CK2), .D(g8780), .SE(SE), .SI(g560), .Q(g617));
S_DFFX1 S_DFF_262 (.CK(CK2), .D(g4894), .SE(SE), .SI(g617), .Q(g17));
S_DFFX1 S_DFF_263 (.CK(CK2), .D(g11653), .SE(SE), .SI(g17), .Q(g336));
S_DFFX1 S_DFF_264 (.CK(CK2), .D(g11466), .SE(SE), .SI(g336), .Q(g456));
S_DFFX1 S_DFF_265 (.CK(CK2), .D(g5643), .SE(SE), .SI(g456), .Q(g305));
S_DFFX1 S_DFF_266 (.CK(CK2), .D(g11642), .SE(SE), .SI(g305), .Q(g345));
S_DFFX1 S_DFF_267 (.CK(CK2), .D(g2613), .SE(SE), .SI(g345), .Q(g8));
S_DFFX1 S_DFF_268 (.CK(CK2), .D(g7811), .SE(SE), .SI(g8), .Q(g1771));
S_DFFX1 S_DFF_269 (.CK(CK2), .D(g8275), .SE(SE), .SI(g1771), .Q(g865));
S_DFFX1 S_DFF_270 (.CK(CK2), .D(g7751), .SE(SE), .SI(g865), .Q(g255));
S_DFFX1 S_DFF_271 (.CK(CK2), .D(g9356), .SE(SE), .SI(g255), .Q(g1945));
S_DFFX1 S_DFF_272 (.CK(CK2), .D(g5661), .SE(SE), .SI(g1945), .Q(g1738));
S_DFFX1 S_DFF_273 (.CK(CK2), .D(g8442), .SE(SE), .SI(g1738), .Q(g1478));
S_DFFX1 S_DFF_274 (.CK(CK2), .D(g7787), .SE(SE), .SI(g1478), .Q(g1035));
S_DFFX1 S_DFF_275 (.CK(CK2), .D(g4217), .SE(SE), .SI(g1035), .Q(g1959));
S_DFFX1 S_DFF_276 (.CK(CK2), .D(g6844), .SE(SE), .SI(g1959), .Q(g1690));
S_DFFX1 S_DFF_277 (.CK(CK2), .D(g8443), .SE(SE), .SI(g1690), .Q(g1482));
S_DFFX1 S_DFF_278 (.CK(CK2), .D(g6817), .SE(SE), .SI(g1482), .Q(g1110));
S_DFFX1 S_DFF_279 (.CK(CK2), .D(g7771), .SE(SE), .SI(g1110), .Q(g296));
S_DFFX1 S_DFF_280 (.CK(CK2), .D(g11034), .SE(SE), .SI(g296), .Q(g1663));
S_DFFX1 S_DFF_281 (.CK(CK2), .D(g8431), .SE(SE), .SI(g1663), .Q(g700));
S_DFFX1 S_DFF_282 (.CK(CK2), .D(g5669), .SE(SE), .SI(g700), .Q(g1762));
S_DFFX1 S_DFF_283 (.CK(CK2), .D(g11510), .SE(SE), .SI(g1762), .Q(g360));
S_DFFX1 S_DFF_284 (.CK(CK2), .D(g6837), .SE(SE), .SI(g360), .Q(g192));
S_DFFX1 S_DFF_285 (.CK(CK2), .D(g10875), .SE(SE), .SI(g192), .Q(g1657));
S_DFFX1 S_DFF_286 (.CK(CK2), .D(g9346), .SE(SE), .SI(g1657), .Q(g722));
S_DFFX1 S_DFF_287 (.CK(CK2), .D(g7780), .SE(SE), .SI(g722), .Q(g61));
S_DFFX1 S_DFF_288 (.CK(CK2), .D(g11051), .SE(SE), .SI(g61), .Q(g566));
S_DFFX1 S_DFF_289 (.CK(CK2), .D(g7809), .SE(SE), .SI(g566), .Q(g1394));
S_DFFX1 S_DFF_290 (.CK(CK2), .D(g6809), .SE(SE), .SI(g1394), .Q(g1089));
S_DFFX1 S_DFF_291 (.CK(CK2), .D(g4897), .SE(SE), .SI(g1089), .Q(g883));
S_DFFX1 S_DFF_292 (.CK(CK2), .D(g6804), .SE(SE), .SI(g883), .Q(g1071));
S_DFFX1 S_DFF_293 (.CK(CK2), .D(g11473), .SE(SE), .SI(g1071), .Q(g986));
S_DFFX1 S_DFF_294 (.CK(CK2), .D(g11470), .SE(SE), .SI(g986), .Q(g971));
S_DFFX1 S_DFF_295 (.CK(CK2), .D(g6338), .SE(SE), .SI(g971), .Q(g1955));
S_DFFX1 S_DFF_296 (.CK(CK2), .D(g7746), .SE(SE), .SI(g1955), .Q(g143));
S_DFFX1 S_DFF_297 (.CK(CK2), .D(g9825), .SE(SE), .SI(g143), .Q(g1814));
S_DFFX1 S_DFF_298 (.CK(CK2), .D(g7797), .SE(SE), .SI(g1814), .Q(g1038));
S_DFFX1 S_DFF_299 (.CK(CK2), .D(g1217), .SE(SE), .SI(g1038), .Q(g1212));
S_DFFX1 S_DFF_300 (.CK(CK2), .D(g9353), .SE(SE), .SI(g1212), .Q(g1918));
S_DFFX1 S_DFF_301 (.CK(CK2), .D(g8273), .SE(SE), .SI(g1918), .Q(g782));
S_DFFX1 S_DFF_302 (.CK(CK2), .D(g9826), .SE(SE), .SI(g782), .Q(g1822));
S_DFFX1 S_DFF_303 (.CK(CK2), .D(g7306), .SE(SE), .SI(g1822), .Q(g237));
S_DFFX1 S_DFF_304 (.CK(CK2), .D(g2638), .SE(SE), .SI(g237), .Q(g746));
S_DFFX1 S_DFF_305 (.CK(CK2), .D(g7795), .SE(SE), .SI(g746), .Q(g1062));
S_DFFX1 S_DFF_306 (.CK(CK2), .D(g8438), .SE(SE), .SI(g1062), .Q(g1462));
S_DFFX1 S_DFF_307 (.CK(CK2), .D(g7748), .SE(SE), .SI(g1462), .Q(g178));
S_DFFX1 S_DFF_308 (.CK(CK2), .D(g11512), .SE(SE), .SI(g178), .Q(g366));
S_DFFX1 S_DFF_309 (.CK(CK2), .D(g4184), .SE(SE), .SI(g366), .Q(g837));
S_DFFX1 S_DFF_310 (.CK(CK2), .D(g9819), .SE(SE), .SI(g837), .Q(g599));
S_DFFX1 S_DFF_311 (.CK(CK2), .D(g11408), .SE(SE), .SI(g599), .Q(g1854));
S_DFFX1 S_DFF_312 (.CK(CK2), .D(g11398), .SE(SE), .SI(g1854), .Q(g944));
S_DFFX1 S_DFF_313 (.CK(CK2), .D(g8287), .SE(SE), .SI(g944), .Q(g1941));
S_DFFX1 S_DFF_314 (.CK(CK2), .D(g8422), .SE(SE), .SI(g1941), .Q(g170));
S_DFFX1 S_DFF_315 (.CK(CK2), .D(g7334), .SE(SE), .SI(g170), .Q(g1520));
S_DFFX1 S_DFF_316 (.CK(CK2), .D(g9342), .SE(SE), .SI(g1520), .Q(g686));
S_DFFX1 S_DFF_317 (.CK(CK2), .D(g11401), .SE(SE), .SI(g686), .Q(g953));
S_DFFX1 S_DFF_318 (.CK(CK2), .D(g6339), .SE(SE), .SI(g953), .Q(g1958));
S_DFFX1 S_DFF_319 (.CK(CK2), .D(g10775), .SE(SE), .SI(g1958), .Q(g40));
S_DFFX1 S_DFF_320 (.CK(CK2), .D(g3329), .SE(SE), .SI(g40), .Q(g1765));
S_DFFX1 S_DFF_321 (.CK(CK2), .D(g10882), .SE(SE), .SI(g1765), .Q(g1733));
S_DFFX1 S_DFF_322 (.CK(CK2), .D(g7303), .SE(SE), .SI(g1733), .Q(g1270));
S_DFFX1 S_DFF_323 (.CK(CK2), .D(g6845), .SE(SE), .SI(g1270), .Q(g1610));
S_DFFX1 S_DFF_324 (.CK(CK2), .D(g8280), .SE(SE), .SI(g1610), .Q(g1796));
S_DFFX1 S_DFF_325 (.CK(CK2), .D(g11632), .SE(SE), .SI(g1796), .Q(g1324));
S_DFFX1 S_DFF_326 (.CK(CK2), .D(g7343), .SE(SE), .SI(g1324), .Q(g1540));
S_DFFX1 S_DFF_327 (.CK(CK2), .D(g7312), .SE(SE), .SI(g1540), .Q(g1377));
S_DFFX1 S_DFF_328 (.CK(CK2), .D(g4898), .SE(SE), .SI(g1377), .Q(g1206));
S_DFFX1 S_DFF_329 (.CK(CK2), .D(g11332), .SE(SE), .SI(g1206), .Q(g491));
S_DFFX1 S_DFF_330 (.CK(CK2), .D(g5670), .SE(SE), .SI(g491), .Q(g1849));
S_DFFX1 S_DFF_331 (.CK(CK2), .D(g7313), .SE(SE), .SI(g1849), .Q(g213));
S_DFFX1 S_DFF_332 (.CK(CK2), .D(g7813), .SE(SE), .SI(g213), .Q(g1781));
S_DFFX1 S_DFF_333 (.CK(CK2), .D(g9351), .SE(SE), .SI(g1781), .Q(g1900));
S_DFFX1 S_DFF_334 (.CK(CK2), .D(g7298), .SE(SE), .SI(g1900), .Q(g1245));
S_DFFX1 S_DFF_335 (.CK(CK2), .D(g11593), .SE(SE), .SI(g1245), .Q(g108));
S_DFFX1 S_DFF_336 (.CK(CK2), .D(g7287), .SE(SE), .SI(g108), .Q(g630));
S_DFFX1 S_DFF_337 (.CK(CK2), .D(g8427), .SE(SE), .SI(g630), .Q(g148));
S_DFFX1 S_DFF_338 (.CK(CK2), .D(g4183), .SE(SE), .SI(g148), .Q(g833));
S_DFFX1 S_DFF_339 (.CK(CK2), .D(g8285), .SE(SE), .SI(g833), .Q(g1923));
S_DFFX1 S_DFF_340 (.CK(CK2), .D(g8571), .SE(SE), .SI(g1923), .Q(g936));
S_DFFX1 S_DFF_341 (.CK(CK2), .D(g6315), .SE(SE), .SI(g936), .Q(g1215));
S_DFFX1 S_DFF_342 (.CK(CK2), .D(g11629), .SE(SE), .SI(g1215), .Q(g1314));
S_DFFX1 S_DFF_343 (.CK(CK2), .D(g4187), .SE(SE), .SI(g1314), .Q(g849));
S_DFFX1 S_DFF_344 (.CK(CK2), .D(g11654), .SE(SE), .SI(g849), .Q(g1336));
S_DFFX1 S_DFF_345 (.CK(CK2), .D(g7763), .SE(SE), .SI(g1336), .Q(g272));
S_DFFX1 S_DFF_346 (.CK(CK2), .D(g8573), .SE(SE), .SI(g272), .Q(g1806));
S_DFFX1 S_DFF_347 (.CK(CK2), .D(g8568), .SE(SE), .SI(g1806), .Q(g826));
S_DFFX1 S_DFF_348 (.CK(CK2), .D(g7796), .SE(SE), .SI(g826), .Q(g1065));
S_DFFX1 S_DFF_349 (.CK(CK2), .D(g8281), .SE(SE), .SI(g1065), .Q(g1887));
S_DFFX1 S_DFF_350 (.CK(CK2), .D(g10871), .SE(SE), .SI(g1887), .Q(g37));
S_DFFX1 S_DFF_351 (.CK(CK2), .D(g11406), .SE(SE), .SI(g37), .Q(g968));
S_DFFX1 S_DFF_352 (.CK(CK2), .D(g5673), .SE(SE), .SI(g968), .Q(g1845));
S_DFFX1 S_DFF_353 (.CK(CK2), .D(g6310), .SE(SE), .SI(g1845), .Q(g1137));
S_DFFX1 S_DFF_354 (.CK(CK2), .D(g9350), .SE(SE), .SI(g1137), .Q(g1891));
S_DFFX1 S_DFF_355 (.CK(CK2), .D(g7300), .SE(SE), .SI(g1891), .Q(g1255));
S_DFFX1 S_DFF_356 (.CK(CK2), .D(g7753), .SE(SE), .SI(g1255), .Q(g257));
S_DFFX1 S_DFF_357 (.CK(CK2), .D(g9821), .SE(SE), .SI(g257), .Q(g874));
S_DFFX1 S_DFF_358 (.CK(CK2), .D(g9818), .SE(SE), .SI(g874), .Q(g591));
S_DFFX1 S_DFF_359 (.CK(CK2), .D(g9347), .SE(SE), .SI(g591), .Q(g731));
S_DFFX1 S_DFF_360 (.CK(CK2), .D(g8781), .SE(SE), .SI(g731), .Q(g636));
S_DFFX1 S_DFF_361 (.CK(CK2), .D(g8276), .SE(SE), .SI(g636), .Q(g1218));
S_DFFX1 S_DFF_362 (.CK(CK2), .D(g9820), .SE(SE), .SI(g1218), .Q(g605));
S_DFFX1 S_DFF_363 (.CK(CK2), .D(g7776), .SE(SE), .SI(g605), .Q(g79));
S_DFFX1 S_DFF_364 (.CK(CK2), .D(g7749), .SE(SE), .SI(g79), .Q(g182));
S_DFFX1 S_DFF_365 (.CK(CK2), .D(g11400), .SE(SE), .SI(g182), .Q(g950));
S_DFFX1 S_DFF_366 (.CK(CK2), .D(g6308), .SE(SE), .SI(g950), .Q(g1129));
S_DFFX1 S_DFF_367 (.CK(CK2), .D(g4189), .SE(SE), .SI(g1129), .Q(g857));
BUFX1 S_BUFX1_SO (.A(g857), .Y(SO));
DFFX1 DFF_368 (.CK(CK1), .D(g11258), .Q(g448));
DFFX1 DFF_369 (.CK(CK1), .D(g9827), .Q(g1828));
DFFX1 DFF_370 (.CK(CK1), .D(g10880), .Q(g1727));
DFFX1 DFF_371 (.CK(CK1), .D(g7360), .Q(g1592));
DFFX1 DFF_372 (.CK(CK1), .D(g6843), .Q(g1703));
DFFX1 DFF_373 (.CK(CK1), .D(g8286), .Q(g1932));
DFFX1 DFF_374 (.CK(CK1), .D(g8870), .Q(g1624));
DFFX1 DFF_375 (.CK(CK1), .D(g4885), .Q(g26));
DFFX1 DFF_376 (.CK(CK1), .D(g6803), .Q(g1068));
DFFX1 DFF_377 (.CK(CK1), .D(g6286), .Q(g578));
DFFX1 DFF_378 (.CK(CK1), .D(g11260), .Q(g440));
DFFX1 DFF_379 (.CK(CK1), .D(g11338), .Q(g476));
DFFX1 DFF_380 (.CK(CK1), .D(g7745), .Q(g119));
DFFX1 DFF_381 (.CK(CK1), .D(g9340), .Q(g668));
DFFX1 DFF_382 (.CK(CK1), .D(g8418), .Q(g139));
DFFX1 DFF_383 (.CK(CK1), .D(g6305), .Q(g1149));
DFFX1 DFF_384 (.CK(CK1), .D(g10868), .Q(g34));
DFFX1 DFF_385 (.CK(CK1), .D(g7366), .Q(g1848));
DFFX1 DFF_386 (.CK(CK1), .D(g7760), .Q(g263));
DFFX1 DFF_387 (.CK(CK1), .D(g8274), .Q(g818));
DFFX1 DFF_388 (.CK(CK1), .D(g5664), .Q(g1747));
DFFX1 DFF_389 (.CK(CK1), .D(g6802), .Q(g802));
DFFX1 DFF_390 (.CK(CK1), .D(g7764), .Q(g275));
DFFX1 DFF_391 (.CK(CK1), .D(g7338), .Q(g1524));
DFFX1 DFF_392 (.CK(CK1), .D(g7355), .Q(g1577));
DFFX1 DFF_393 (.CK(CK1), .D(g7786), .Q(g810));
DFFX1 DFF_394 (.CK(CK1), .D(g11264), .Q(g391));
DFFX1 DFF_395 (.CK(CK1), .D(g9339), .Q(g658));
DFFX1 DFF_396 (.CK(CK1), .D(g7318), .Q(g1386));
DFFX1 DFF_397 (.CK(CK1), .D(g7750), .Q(g253));
DFFX1 DFF_398 (.CK(CK1), .D(g9822), .Q(g875));
DFFX1 DFF_399 (.CK(CK1), .D(g6307), .Q(g1125));
DFFX1 DFF_400 (.CK(CK1), .D(g7304), .Q(g201));
DFFX1 DFF_401 (.CK(CK1), .D(g7295), .Q(g1280));
DFFX1 DFF_402 (.CK(CK1), .D(g6807), .Q(g1083));
DFFX1 DFF_403 (.CK(CK1), .D(g8066), .Q(g650));
DFFX1 DFF_404 (.CK(CK1), .D(g8874), .Q(g1636));
DFFX1 DFF_405 (.CK(CK1), .D(g4188), .Q(g853));
DFFX1 DFF_406 (.CK(CK1), .D(g11270), .Q(g421));
DFFX1 DFF_407 (.CK(CK1), .D(g6798), .Q(g762));
DFFX1 DFF_408 (.CK(CK1), .D(g11402), .Q(g956));
DFFX1 DFF_409 (.CK(CK1), .D(g11441), .Q(g378));
DFFX1 DFF_410 (.CK(CK1), .D(g5667), .Q(g1756));
DFFX1 DFF_411 (.CK(CK1), .D(g6297), .Q(g589));
DFFX1 DFF_412 (.CK(CK1), .D(g4185), .Q(g841));
DFFX1 DFF_413 (.CK(CK1), .D(g7798), .Q(g1027));
DFFX1 DFF_414 (.CK(CK1), .D(g7803), .Q(g1003));
DFFX1 DFF_415 (.CK(CK1), .D(g8991), .Q(g1403));
DFFX1 DFF_416 (.CK(CK1), .D(g6312), .Q(g1145));
DFFX1 DFF_417 (.CK(CK1), .D(g6816), .Q(g1107));
DFFX1 DFF_418 (.CK(CK1), .D(g8277), .Q(g1223));
DFFX1 DFF_419 (.CK(CK1), .D(g11267), .Q(g406));
DFFX1 DFF_420 (.CK(CK1), .D(g11185), .Q(g1811));
DFFX1 DFF_421 (.CK(CK1), .D(g11183), .Q(g1642));
DFFX1 DFF_422 (.CK(CK1), .D(g7790), .Q(g1047));
DFFX1 DFF_423 (.CK(CK1), .D(g10874), .Q(g1654));
DFFX1 DFF_424 (.CK(CK1), .D(g6835), .Q(g197));
DFFX1 DFF_425 (.CK(CK1), .D(g7361), .Q(g1595));
DFFX1 DFF_426 (.CK(CK1), .D(g7342), .Q(g1537));
DFFX1 DFF_427 (.CK(CK1), .D(g8434), .Q(g727));
DFFX1 DFF_428 (.CK(CK1), .D(g7804), .Q(g999));
DFFX1 DFF_429 (.CK(CK1), .D(g6801), .Q(g798));
DFFX1 DFF_430 (.CK(CK1), .D(g11324), .Q(g481));
DFFX1 DFF_431 (.CK(CK1), .D(g4895), .Q(g754));
DFFX1 DFF_432 (.CK(CK1), .D(g11634), .Q(g1330));
DFFX1 DFF_433 (.CK(CK1), .D(g4186), .Q(g845));
DFFX1 DFF_434 (.CK(CK1), .D(g8567), .Q(g790));
DFFX1 DFF_435 (.CK(CK1), .D(g8449), .Q(g1512));
DFFX1 DFF_436 (.CK(CK1), .D(g113), .Q(g114));
DFFX1 DFF_437 (.CK(CK1), .D(g8445), .Q(g1490));
DFFX1 DFF_438 (.CK(CK1), .D(g6300), .Q(g1166));
DFFX1 DFF_439 (.CK(CK1), .D(g7793), .Q(g1056));
DFFX1 DFF_440 (.CK(CK1), .D(g11506), .Q(g348));
DFFX1 DFF_441 (.CK(CK1), .D(g874), .Q(g868));
DFFX1 DFF_442 (.CK(CK1), .D(g7301), .Q(g1260));
DFFX1 DFF_443 (.CK(CK1), .D(g7756), .Q(g260));
DFFX1 DFF_444 (.CK(CK1), .D(g8420), .Q(g131));
DFFX1 DFF_445 (.CK(CK1), .D(g2731), .Q(g7));
DFFX1 DFF_446 (.CK(CK1), .D(g7754), .Q(g258));
DFFX1 DFF_447 (.CK(CK1), .D(g11330), .Q(g521));
DFFX1 DFF_448 (.CK(CK1), .D(g11630), .Q(g1318));
DFFX1 DFF_449 (.CK(CK1), .D(g9348), .Q(g1872));
DFFX1 DFF_450 (.CK(CK1), .D(g9341), .Q(g677));
DFFX1 DFF_451 (.CK(CK1), .D(g6290), .Q(g582));
DFFX1 DFF_452 (.CK(CK1), .D(g7320), .Q(g1393));
DFFX1 DFF_453 (.CK(CK1), .D(g7346), .Q(g1549));
DFFX1 DFF_454 (.CK(CK1), .D(g11399), .Q(g947));
DFFX1 DFF_455 (.CK(CK1), .D(g9895), .Q(g1834));
DFFX1 DFF_456 (.CK(CK1), .D(g7362), .Q(g1598));
DFFX1 DFF_457 (.CK(CK1), .D(g6306), .Q(g1121));
DFFX1 DFF_458 (.CK(CK1), .D(g11631), .Q(g1321));
DFFX1 DFF_459 (.CK(CK1), .D(g11335), .Q(g506));
DFFX1 DFF_460 (.CK(CK1), .D(g11043), .Q(g546));
DFFX1 DFF_461 (.CK(CK1), .D(g9352), .Q(g1909));
DFFX1 DFF_462 (.CK(CK1), .D(g6298), .Q(g755));
DFFX1 DFF_463 (.CK(CK1), .D(g7347), .Q(g1552));
DFFX1 DFF_464 (.CK(CK1), .D(g6292), .Q(g584));
DFFX1 DFF_465 (.CK(CK1), .D(g11042), .Q(g1687));
DFFX1 DFF_466 (.CK(CK1), .D(g7358), .Q(g1586));
DFFX1 DFF_467 (.CK(CK1), .D(g5648), .Q(g324));
DFFX1 DFF_468 (.CK(CK1), .D(g6311), .Q(g1141));
DFFX1 DFF_469 (.CK(CK1), .D(g4900), .Q(g1570));
DFFX1 DFF_470 (.CK(CK1), .D(g11655), .Q(g1341));
DFFX1 DFF_471 (.CK(CK1), .D(g4901), .Q(g1710));
DFFX1 DFF_472 (.CK(CK1), .D(g11184), .Q(g1645));
DFFX1 DFF_473 (.CK(CK1), .D(g7321), .Q(g115));
DFFX1 DFF_474 (.CK(CK1), .D(g8419), .Q(g135));
DFFX1 DFF_475 (.CK(CK1), .D(g11329), .Q(g525));
DFFX1 DFF_476 (.CK(CK1), .D(g6289), .Q(g581));
DFFX1 DFF_477 (.CK(CK1), .D(g7365), .Q(g1607));
DFFX1 DFF_478 (.CK(CK1), .D(g5647), .Q(g321));
DFFX1 DFF_479 (.CK(CK1), .D(g7782), .Q(g67));
DFFX1 DFF_480 (.CK(CK1), .D(g11443), .Q(g1275));
DFFX1 DFF_481 (.CK(CK1), .D(g11628), .Q(g1311));
DFFX1 DFF_482 (.CK(CK1), .D(g8868), .Q(g1615));
DFFX1 DFF_483 (.CK(CK1), .D(g11442), .Q(g382));
DFFX1 DFF_484 (.CK(CK1), .D(g6825), .Q(g1374));
DFFX1 DFF_485 (.CK(CK1), .D(g7761), .Q(g266));
DFFX1 DFF_486 (.CK(CK1), .D(g7294), .Q(g1284));
DFFX1 DFF_487 (.CK(CK1), .D(g7314), .Q(g1380));
DFFX1 DFF_488 (.CK(CK1), .D(g8428), .Q(g673));
DFFX1 DFF_489 (.CK(CK1), .D(g5672), .Q(g1853));
DFFX1 DFF_490 (.CK(CK1), .D(g8424), .Q(g162));
DFFX1 DFF_491 (.CK(CK1), .D(g11268), .Q(g411));
DFFX1 DFF_492 (.CK(CK1), .D(g11262), .Q(g431));
DFFX1 DFF_493 (.CK(CK1), .D(g8283), .Q(g1905));
DFFX1 DFF_494 (.CK(CK1), .D(g7333), .Q(g1515));
DFFX1 DFF_495 (.CK(CK1), .D(g8872), .Q(g1630));
DFFX1 DFF_496 (.CK(CK1), .D(g7774), .Q(g49));
DFFX1 DFF_497 (.CK(CK1), .D(g7802), .Q(g991));
DFFX1 DFF_498 (.CK(CK1), .D(g7291), .Q(g1300));
DFFX1 DFF_499 (.CK(CK1), .D(g11505), .Q(g339));
DFFX1 DFF_500 (.CK(CK1), .D(g7752), .Q(g256));
DFFX1 DFF_501 (.CK(CK1), .D(g5665), .Q(g1750));
DFFX1 DFF_502 (.CK(CK1), .D(g6293), .Q(g585));
DFFX1 DFF_503 (.CK(CK1), .D(g8988), .Q(g1440));
DFFX1 DFF_504 (.CK(CK1), .D(g11035), .Q(g1666));
DFFX1 DFF_505 (.CK(CK1), .D(g7339), .Q(g1528));
DFFX1 DFF_506 (.CK(CK1), .D(g11657), .Q(g1351));
DFFX1 DFF_507 (.CK(CK1), .D(g11181), .Q(g1648));
DFFX1 DFF_508 (.CK(CK1), .D(g8421), .Q(g127));
DFFX1 DFF_509 (.CK(CK1), .D(g11611), .Q(g1618));
DFFX1 DFF_510 (.CK(CK1), .D(g7296), .Q(g1235));
DFFX1 DFF_511 (.CK(CK1), .D(g7772), .Q(g299));
DFFX1 DFF_512 (.CK(CK1), .D(g11261), .Q(g435));
DFFX1 DFF_513 (.CK(CK1), .D(g7781), .Q(g64));
DFFX1 DFF_514 (.CK(CK1), .D(g7348), .Q(g1555));
DFFX1 DFF_515 (.CK(CK1), .D(g7801), .Q(g995));
DFFX1 DFF_516 (.CK(CK1), .D(g8869), .Q(g1621));
DFFX1 DFF_517 (.CK(CK1), .D(g6313), .Q(g1113));
DFFX1 DFF_518 (.CK(CK1), .D(g8064), .Q(g643));
DFFX1 DFF_519 (.CK(CK1), .D(g8446), .Q(g1494));
DFFX1 DFF_520 (.CK(CK1), .D(g7352), .Q(g1567));
DFFX1 DFF_521 (.CK(CK1), .D(g8430), .Q(g691));
DFFX1 DFF_522 (.CK(CK1), .D(g11327), .Q(g534));
DFFX1 DFF_523 (.CK(CK1), .D(g7812), .Q(g1776));
DFFX1 DFF_524 (.CK(CK1), .D(g10876), .Q(g569));
DFFX1 DFF_525 (.CK(CK1), .D(g6302), .Q(g1160));
DFFX1 DFF_526 (.CK(CK1), .D(g9824), .Q(g1360));
DFFX1 DFF_527 (.CK(CK1), .D(g7791), .Q(g1050));
DFFX1 DFF_528 (.CK(CK1), .D(g8078), .Q(g1));
DFFX1 DFF_529 (.CK(CK1), .D(g11336), .Q(g511));
DFFX1 DFF_530 (.CK(CK1), .D(g10879), .Q(g1724));
DFFX1 DFF_531 (.CK(CK1), .D(g7337), .Q(g12));
DFFX1 DFF_532 (.CK(CK1), .D(g8695), .Q(g1878));
DFFX1 DFF_533 (.CK(CK1), .D(g7784), .Q(g73));
INVX1 NOT_0 (.Y(I8854),.A(g4500));
INVX1 NOT_1 (.Y(g5652),.A(I9117));
INVX1 NOT_2 (.Y(I12913),.A(g7845));
INVX1 NOT_3 (.Y(g11354),.A(I17179));
INVX1 NOT_4 (.Y(g6837),.A(I10891));
INVX1 NOT_5 (.Y(I10941),.A(g6555));
INVX1 NOT_6 (.Y(I6979),.A(g2888));
INVX1 NOT_7 (.Y(g5843),.A(I9458));
INVX1 NOT_8 (.Y(g2771),.A(I5854));
INVX1 NOT_9 (.Y(g3537),.A(g3164));
INVX1 NOT_10 (.Y(g6062),.A(I9699));
INVX1 NOT_11 (.Y(I9984),.A(g5529));
INVX1 NOT_12 (.Y(I14382),.A(g8886));
INVX1 NOT_13 (.Y(g7706),.A(I12335));
INVX1 NOT_14 (.Y(I13618),.A(g8345));
INVX1 NOT_15 (.Y(I15181),.A(g9968));
INVX1 NOT_16 (.Y(g6620),.A(I10573));
INVX1 NOT_17 (.Y(I12436),.A(g7659));
INVX1 NOT_18 (.Y(g5193),.A(g4682));
INVX1 NOT_19 (.Y(g6462),.A(I10394));
INVX1 NOT_20 (.Y(g8925),.A(I14252));
INVX1 NOT_21 (.Y(I14519),.A(g9106));
INVX1 NOT_22 (.Y(g10289),.A(I15691));
INVX1 NOT_23 (.Y(I14176),.A(g8784));
INVX1 NOT_24 (.Y(I14185),.A(g8790));
INVX1 NOT_25 (.Y(g11181),.A(I16944));
INVX1 NOT_26 (.Y(I14675),.A(g9263));
INVX1 NOT_27 (.Y(g2299),.A(g1707));
INVX1 NOT_28 (.Y(I12607),.A(g7633));
INVX1 NOT_29 (.Y(g3272),.A(g2450));
INVX1 NOT_30 (.Y(g2547),.A(g23));
INVX1 NOT_31 (.Y(g9291),.A(g8892));
INVX1 NOT_32 (.Y(I6001),.A(g2548));
INVX1 NOT_33 (.Y(I7048),.A(g2807));
INVX1 NOT_34 (.Y(g10309),.A(I15733));
INVX1 NOT_35 (.Y(g7029),.A(I11180));
INVX1 NOT_36 (.Y(g4440),.A(g4130));
INVX1 NOT_37 (.Y(I9544),.A(g5024));
INVX1 NOT_38 (.Y(g10288),.A(I15688));
INVX1 NOT_39 (.Y(I12274),.A(g7110));
INVX1 NOT_40 (.Y(I9483),.A(g5050));
INVX1 NOT_41 (.Y(g7787),.A(I12526));
INVX1 NOT_42 (.Y(I6676),.A(g2759));
INVX1 NOT_43 (.Y(I8520),.A(g4338));
INVX1 NOT_44 (.Y(g10571),.A(I16236));
INVX1 NOT_45 (.Y(I17692),.A(g11596));
INVX1 NOT_46 (.Y(I17761),.A(g11652));
INVX1 NOT_47 (.Y(I13469),.A(g8147));
INVX1 NOT_48 (.Y(g9344),.A(I14537));
INVX1 NOT_49 (.Y(g7956),.A(g7432));
INVX1 NOT_50 (.Y(g3417),.A(I6624));
INVX1 NOT_51 (.Y(g4323),.A(g4130));
INVX1 NOT_52 (.Y(I11286),.A(g6551));
INVX1 NOT_53 (.Y(I8031),.A(g3540));
INVX1 NOT_54 (.Y(g7675),.A(I12300));
INVX1 NOT_55 (.Y(g8320),.A(I13344));
INVX1 NOT_56 (.Y(I12565),.A(g7388));
INVX1 NOT_57 (.Y(I16644),.A(g10865));
INVX1 NOT_58 (.Y(I11306),.A(g6731));
INVX1 NOT_59 (.Y(g1981),.A(g650));
INVX1 NOT_60 (.Y(I7333),.A(g3729));
INVX1 NOT_61 (.Y(I13039),.A(g8054));
INVX1 NOT_62 (.Y(g3982),.A(g3052));
INVX1 NOT_63 (.Y(g6249),.A(I10006));
INVX1 NOT_64 (.Y(g9259),.A(g8892));
INVX1 NOT_65 (.Y(I15190),.A(g9974));
INVX1 NOT_66 (.Y(g11426),.A(I17331));
INVX1 NOT_67 (.Y(g9819),.A(I14958));
INVX1 NOT_68 (.Y(g8277),.A(I13203));
INVX1 NOT_69 (.Y(I5050),.A(g1216));
INVX1 NOT_70 (.Y(I5641),.A(g546));
INVX1 NOT_71 (.Y(g5121),.A(g4682));
INVX1 NOT_72 (.Y(g1997),.A(g798));
INVX1 NOT_73 (.Y(g3629),.A(g3228));
INVX1 NOT_74 (.Y(g3328),.A(I6501));
INVX1 NOT_75 (.Y(I12641),.A(g7709));
INVX1 NOT_76 (.Y(g5670),.A(I9171));
INVX1 NOT_77 (.Y(g6842),.A(I10898));
INVX1 NOT_78 (.Y(g8617),.A(g8465));
INVX1 NOT_79 (.Y(I15520),.A(g10035));
INVX1 NOT_80 (.Y(I7396),.A(g4102));
INVX1 NOT_81 (.Y(I7803),.A(g3820));
INVX1 NOT_82 (.Y(g3330),.A(I6507));
INVX1 NOT_83 (.Y(g2991),.A(I6233));
INVX1 NOT_84 (.Y(I9461),.A(g4940));
INVX1 NOT_85 (.Y(g2244),.A(I5251));
INVX1 NOT_86 (.Y(g6192),.A(I9923));
INVX1 NOT_87 (.Y(g6298),.A(I10153));
INVX1 NOT_88 (.Y(g6085),.A(I9734));
INVX1 NOT_89 (.Y(I12153),.A(g6874));
INVX1 NOT_90 (.Y(g4351),.A(I7630));
INVX1 NOT_91 (.Y(I11677),.A(g7056));
INVX1 NOT_92 (.Y(g10687),.A(I16356));
INVX1 NOT_93 (.Y(g4530),.A(I7935));
INVX1 NOT_94 (.Y(g8516),.A(I13717));
INVX1 NOT_95 (.Y(g5232),.A(g4640));
INVX1 NOT_96 (.Y(I13975),.A(g8588));
INVX1 NOT_97 (.Y(g2078),.A(g135));
INVX1 NOT_98 (.Y(I8911),.A(g4565));
INVX1 NOT_99 (.Y(g2340),.A(g1918));
INVX1 NOT_100 (.Y(g7684),.A(g7148));
INVX1 NOT_101 (.Y(I12409),.A(g7501));
INVX1 NOT_102 (.Y(g7745),.A(I12400));
INVX1 NOT_103 (.Y(g8987),.A(I14382));
INVX1 NOT_104 (.Y(g11546),.A(g11519));
INVX1 NOT_105 (.Y(I10729),.A(g5935));
INVX1 NOT_106 (.Y(g5253),.A(g4346));
INVX1 NOT_107 (.Y(g7338),.A(I11662));
INVX1 NOT_108 (.Y(I7509),.A(g3566));
INVX1 NOT_109 (.Y(I9427),.A(g4963));
INVX1 NOT_110 (.Y(g3800),.A(g3292));
INVX1 NOT_111 (.Y(I15088),.A(g9832));
INVX1 NOT_112 (.Y(g2907),.A(I6074));
INVX1 NOT_113 (.Y(g7791),.A(I12538));
INVX1 NOT_114 (.Y(I11143),.A(g6446));
INVX1 NOT_115 (.Y(g6854),.A(I10920));
INVX1 NOT_116 (.Y(g11088),.A(I16871));
INVX1 NOT_117 (.Y(g7309),.A(I11575));
INVX1 NOT_118 (.Y(g8299),.A(I13255));
INVX1 NOT_119 (.Y(I9046),.A(g4736));
INVX1 NOT_120 (.Y(g6941),.A(g6503));
INVX1 NOT_121 (.Y(g2435),.A(g201));
INVX1 NOT_122 (.Y(I14439),.A(g8969));
INVX1 NOT_123 (.Y(g4010),.A(g3144));
INVX1 NOT_124 (.Y(g2082),.A(g1371));
INVX1 NOT_125 (.Y(I6932),.A(g2850));
INVX1 NOT_126 (.Y(I7662),.A(g3336));
INVX1 NOT_127 (.Y(I9446),.A(g5052));
INVX1 NOT_128 (.Y(g5519),.A(g4811));
INVX1 NOT_129 (.Y(g5740),.A(I9302));
INVX1 NOT_130 (.Y(I5289),.A(g49));
INVX1 NOT_131 (.Y(I9514),.A(g5094));
INVX1 NOT_132 (.Y(g7808),.A(I12589));
INVX1 NOT_133 (.Y(g2482),.A(I5565));
INVX1 NOT_134 (.Y(I5658),.A(g560));
INVX1 NOT_135 (.Y(I15497),.A(g10119));
INVX1 NOT_136 (.Y(I6624),.A(g2629));
INVX1 NOT_137 (.Y(g8892),.A(I14242));
INVX1 NOT_138 (.Y(I11169),.A(g6481));
INVX1 NOT_139 (.Y(g3213),.A(I6388));
INVX1 NOT_140 (.Y(I6068),.A(g2227));
INVX1 NOT_141 (.Y(g11497),.A(I17510));
INVX1 NOT_142 (.Y(I13791),.A(g8518));
INVX1 NOT_143 (.Y(I16867),.A(g10913));
INVX1 NOT_144 (.Y(I10349),.A(g6215));
INVX1 NOT_145 (.Y(g10260),.A(g10125));
INVX1 NOT_146 (.Y(g7759),.A(I12442));
INVX1 NOT_147 (.Y(I8473),.A(g4577));
INVX1 NOT_148 (.Y(I14349),.A(g8958));
INVX1 NOT_149 (.Y(g6708),.A(I10689));
INVX1 NOT_150 (.Y(g10668),.A(g10563));
INVX1 NOT_151 (.Y(I5271),.A(g70));
INVX1 NOT_152 (.Y(I9191),.A(g5546));
INVX1 NOT_153 (.Y(I9391),.A(g5013));
INVX1 NOT_154 (.Y(g6219),.A(g5426));
INVX1 NOT_155 (.Y(I15250),.A(g9980));
INVX1 NOT_156 (.Y(I17100),.A(g11221));
INVX1 NOT_157 (.Y(I14906),.A(g9508));
INVX1 NOT_158 (.Y(g9825),.A(I14976));
INVX1 NOT_159 (.Y(g7201),.A(I11427));
INVX1 NOT_160 (.Y(I14083),.A(g8747));
INVX1 NOT_161 (.Y(g10195),.A(I15559));
INVX1 NOT_162 (.Y(I8324),.A(g4794));
INVX1 NOT_163 (.Y(g6031),.A(I9642));
INVX1 NOT_164 (.Y(g2915),.A(I6094));
INVX1 NOT_165 (.Y(I13666),.A(g8292));
INVX1 NOT_166 (.Y(I9695),.A(g5212));
INVX1 NOT_167 (.Y(I11363),.A(g6595));
INVX1 NOT_168 (.Y(I11217),.A(g6529));
INVX1 NOT_169 (.Y(g6431),.A(g6145));
INVX1 NOT_170 (.Y(g6252),.A(I10015));
INVX1 NOT_171 (.Y(g4172),.A(I7333));
INVX1 NOT_172 (.Y(g6812),.A(I10846));
INVX1 NOT_173 (.Y(g8991),.A(I14394));
INVX1 NOT_174 (.Y(g4372),.A(I7677));
INVX1 NOT_175 (.Y(g7049),.A(I11228));
INVX1 NOT_176 (.Y(I6576),.A(g2617));
INVX1 NOT_177 (.Y(g10525),.A(g10499));
INVX1 NOT_178 (.Y(g10488),.A(I16101));
INVX1 NOT_179 (.Y(I10566),.A(g5904));
INVX1 NOT_180 (.Y(I13478),.A(g8191));
INVX1 NOT_181 (.Y(g5586),.A(I8996));
INVX1 NOT_182 (.Y(g8709),.A(g8674));
INVX1 NOT_183 (.Y(g2214),.A(g115));
INVX1 NOT_184 (.Y(I9536),.A(g5008));
INVX1 NOT_185 (.Y(g6176),.A(I9905));
INVX1 NOT_186 (.Y(g4618),.A(g3829));
INVX1 NOT_187 (.Y(I15296),.A(g9995));
INVX1 NOT_188 (.Y(g4143),.A(I7291));
INVX1 NOT_189 (.Y(I7381),.A(g4078));
INVX1 NOT_190 (.Y(I9159),.A(g5033));
INVX1 NOT_191 (.Y(g11339),.A(I17142));
INVX1 NOT_192 (.Y(g8140),.A(I13017));
INVX1 NOT_193 (.Y(I16979),.A(g11088));
INVX1 NOT_194 (.Y(I16496),.A(g10707));
INVX1 NOT_195 (.Y(g8078),.A(I12936));
INVX1 NOT_196 (.Y(I7847),.A(g3435));
INVX1 NOT_197 (.Y(I9359),.A(g5576));
INVX1 NOT_198 (.Y(g8340),.A(I13400));
INVX1 NOT_199 (.Y(g2110),.A(I5002));
INVX1 NOT_200 (.Y(I15338),.A(g10013));
INVX1 NOT_201 (.Y(g6405),.A(g6133));
INVX1 NOT_202 (.Y(g8478),.A(I13678));
INVX1 NOT_203 (.Y(I16111),.A(g10385));
INVX1 NOT_204 (.Y(g4282),.A(g4013));
INVX1 NOT_205 (.Y(g11644),.A(I17736));
INVX1 NOT_206 (.Y(g7604),.A(I12162));
INVX1 NOT_207 (.Y(g9768),.A(g9432));
INVX1 NOT_208 (.Y(g4566),.A(g3753));
INVX1 NOT_209 (.Y(g7098),.A(I11333));
INVX1 NOT_210 (.Y(g10893),.A(I16641));
INVX1 NOT_211 (.Y(I4961),.A(g254));
INVX1 NOT_212 (.Y(g4988),.A(I8358));
INVX1 NOT_213 (.Y(g6286),.A(I10117));
INVX1 NOT_214 (.Y(g8959),.A(I14326));
INVX1 NOT_215 (.Y(I13580),.A(g8338));
INVX1 NOT_216 (.Y(I9016),.A(g4722));
INVX1 NOT_217 (.Y(I6398),.A(g2335));
INVX1 NOT_218 (.Y(g8517),.A(I13720));
INVX1 NOT_219 (.Y(g3348),.A(g2733));
INVX1 NOT_220 (.Y(I15060),.A(g9696));
INVX1 NOT_221 (.Y(I15968),.A(g10408));
INVX1 NOT_222 (.Y(I5332),.A(g756));
INVX1 NOT_223 (.Y(g8482),.A(g8329));
INVX1 NOT_224 (.Y(g2002),.A(g818));
INVX1 NOT_225 (.Y(I10138),.A(g5677));
INVX1 NOT_226 (.Y(g11060),.A(g10937));
INVX1 NOT_227 (.Y(I17407),.A(g11417));
INVX1 NOT_228 (.Y(I12303),.A(g7242));
INVX1 NOT_229 (.Y(g5645),.A(I9096));
INVX1 NOT_230 (.Y(I15855),.A(g10336));
INVX1 NOT_231 (.Y(g2824),.A(I5932));
INVX1 NOT_232 (.Y(g11197),.A(g11112));
INVX1 NOT_233 (.Y(g4555),.A(I7964));
INVX1 NOT_234 (.Y(g5691),.A(g5236));
INVX1 NOT_235 (.Y(I9642),.A(g5229));
INVX1 NOT_236 (.Y(g7539),.A(I11953));
INVX1 NOT_237 (.Y(g7896),.A(I12678));
INVX1 NOT_238 (.Y(g8656),.A(I13941));
INVX1 NOT_239 (.Y(g9887),.A(I15068));
INVX1 NOT_240 (.Y(I8199),.A(g4013));
INVX1 NOT_241 (.Y(g6974),.A(g6365));
INVX1 NOT_242 (.Y(g6270),.A(I10069));
INVX1 NOT_243 (.Y(I14415),.A(g8940));
INVX1 NOT_244 (.Y(g3260),.A(I6428));
INVX1 NOT_245 (.Y(g11411),.A(I17274));
INVX1 NOT_246 (.Y(I10852),.A(g6751));
INVX1 NOT_247 (.Y(g10042),.A(I15253));
INVX1 NOT_248 (.Y(g10255),.A(g10139));
INVX1 NOT_249 (.Y(g6073),.A(I9712));
INVX1 NOT_250 (.Y(g10189),.A(I15545));
INVX1 NOT_251 (.Y(I4903),.A(g259));
INVX1 NOT_252 (.Y(g2877),.A(I6025));
INVX1 NOT_253 (.Y(I11531),.A(g7126));
INVX1 NOT_254 (.Y(g10679),.A(g10584));
INVX1 NOT_255 (.Y(g6796),.A(g6252));
INVX1 NOT_256 (.Y(I8900),.A(g4560));
INVX1 NOT_257 (.Y(I16735),.A(g10855));
INVX1 NOT_258 (.Y(g1968),.A(g369));
INVX1 NOT_259 (.Y(g5879),.A(I9498));
INVX1 NOT_260 (.Y(I10963),.A(g6793));
INVX1 NOT_261 (.Y(g10270),.A(g10156));
INVX1 NOT_262 (.Y(g3463),.A(g3256));
INVX1 NOT_263 (.Y(g7268),.A(I11505));
INVX1 NOT_264 (.Y(g7362),.A(I11734));
INVX1 NOT_265 (.Y(I11740),.A(g7030));
INVX1 NOT_266 (.Y(g10188),.A(I15542));
INVX1 NOT_267 (.Y(I12174),.A(g6939));
INVX1 NOT_268 (.Y(I12796),.A(g7543));
INVX1 NOT_269 (.Y(g5659),.A(I9138));
INVX1 NOT_270 (.Y(g7419),.A(g7206));
INVX1 NOT_271 (.Y(I15503),.A(g10044));
INVX1 NOT_272 (.Y(I17441),.A(g11445));
INVX1 NOT_273 (.Y(g6980),.A(I11127));
INVX1 NOT_274 (.Y(I17206),.A(g11323));
INVX1 NOT_275 (.Y(g4113),.A(I7255));
INVX1 NOT_276 (.Y(g6069),.A(I9706));
INVX1 NOT_277 (.Y(g11503),.A(I17528));
INVX1 NOT_278 (.Y(g7052),.A(I11235));
INVX1 NOT_279 (.Y(g8110),.A(g7996));
INVX1 NOT_280 (.Y(g2556),.A(g186));
INVX1 NOT_281 (.Y(g4313),.A(g3586));
INVX1 NOT_282 (.Y(I16196),.A(g10496));
INVX1 NOT_283 (.Y(I7817),.A(g3399));
INVX1 NOT_284 (.Y(g8310),.A(I13314));
INVX1 NOT_285 (.Y(g10460),.A(I15971));
INVX1 NOT_286 (.Y(g2222),.A(g158));
INVX1 NOT_287 (.Y(I11953),.A(g6907));
INVX1 NOT_288 (.Y(I13373),.A(g8226));
INVX1 NOT_289 (.Y(I6818),.A(g2758));
INVX1 NOT_290 (.Y(g4202),.A(I7423));
INVX1 NOT_291 (.Y(I6867),.A(g2949));
INVX1 NOT_292 (.Y(I9880),.A(g5405));
INVX1 NOT_293 (.Y(g10093),.A(I15326));
INVX1 NOT_294 (.Y(I10484),.A(g6155));
INVX1 NOT_295 (.Y(g9845),.A(g9679));
INVX1 NOT_296 (.Y(g3720),.A(I6888));
INVX1 NOT_297 (.Y(g10267),.A(g10130));
INVX1 NOT_298 (.Y(g10294),.A(I15704));
INVX1 NOT_299 (.Y(I11800),.A(g7246));
INVX1 NOT_300 (.Y(g4908),.A(g4396));
INVX1 NOT_301 (.Y(g5111),.A(I8499));
INVX1 NOT_302 (.Y(g11450),.A(I17407));
INVX1 NOT_303 (.Y(I13800),.A(g8500));
INVX1 NOT_304 (.Y(g5275),.A(g4371));
DFFX1 DFF_0 (.CK(CK1), .D(g5660), .Q(g1289));
DFFX1 DFF_1 (.CK(CK1), .D(g9349), .Q(g1882));
DFFX1 DFF_2 (.CK(CK1), .D(g5644), .Q(g312));
DFFX1 DFF_3 (.CK(CK1), .D(g11257), .Q(g452));
DFFX1 DFF_4 (.CK(CK1), .D(g8272), .Q(g123));
DFFX1 DFF_5 (.CK(CK1), .D(g7315), .Q(g207));
DFFX1 DFF_6 (.CK(CK1), .D(g9345), .Q(g713));
DFFX1 DFF_7 (.CK(CK1), .D(g6304), .Q(g1153));
DFFX1 DFF_8 (.CK(CK1), .D(g10873), .Q(g1209));
DFFX1 DFF_9 (.CK(CK1), .D(g5663), .Q(g1744));
DFFX1 DFF_10 (.CK(CK1), .D(g7349), .Q(g1558));
DFFX1 DFF_11 (.CK(CK1), .D(g9343), .Q(g695));
DFFX1 DFF_12 (.CK(CK1), .D(g11467), .Q(g461));
DFFX1 DFF_13 (.CK(CK1), .D(g8572), .Q(g940));
DFFX1 DFF_14 (.CK(CK1), .D(g11471), .Q(g976));
DFFX1 DFF_15 (.CK(CK1), .D(g8432), .Q(g709));
DFFX1 DFF_16 (.CK(CK1), .D(g6810), .Q(g1092));
INVX1 NOT_305 (.Y(I11417),.A(g6638));
INVX1 NOT_306 (.Y(I17758),.A(g11647));
INVX1 NOT_307 (.Y(g3318),.A(g2245));
INVX1 NOT_308 (.Y(g11315),.A(I17108));
INVX1 NOT_309 (.Y(g4094),.A(g2744));
INVX1 NOT_310 (.Y(I17435),.A(g11454));
INVX1 NOT_311 (.Y(g10065),.A(I15293));
INVX1 NOT_312 (.Y(I5092),.A(g32));
INVX1 NOT_313 (.Y(g8002),.A(I12832));
INVX1 NOT_314 (.Y(g5615),.A(I9043));
INVX1 NOT_315 (.Y(g4567),.A(g3374));
INVX1 NOT_316 (.Y(I8259),.A(g4590));
INVX1 NOT_317 (.Y(g11202),.A(g11112));
INVX1 NOT_318 (.Y(g7728),.A(I12369));
INVX1 NOT_319 (.Y(g6287),.A(I10120));
INVX1 NOT_320 (.Y(I14312),.A(g8814));
INVX1 NOT_321 (.Y(I9612),.A(g5149));
INVX1 NOT_322 (.Y(g10875),.A(I16595));
INVX1 NOT_323 (.Y(I9243),.A(g5245));
INVX1 NOT_324 (.Y(g11055),.A(g10950));
INVX1 NOT_325 (.Y(g3393),.A(g3144));
INVX1 NOT_326 (.Y(g9807),.A(g9490));
INVX1 NOT_327 (.Y(g11111),.A(g10974));
INVX1 NOT_328 (.Y(g4776),.A(g3586));
INVX1 NOT_329 (.Y(I9935),.A(g5477));
INVX1 NOT_330 (.Y(g4593),.A(I8004));
INVX1 NOT_331 (.Y(I11964),.A(g6910));
INVX1 NOT_332 (.Y(I7441),.A(g3473));
INVX1 NOT_333 (.Y(I15986),.A(g10417));
INVX1 NOT_334 (.Y(g3971),.A(I7104));
INVX1 NOT_335 (.Y(g7070),.A(I11289));
INVX1 NOT_336 (.Y(g2237),.A(g713));
INVX1 NOT_337 (.Y(g6399),.A(I10305));
INVX1 NOT_338 (.Y(g5284),.A(g4376));
INVX1 NOT_339 (.Y(I11423),.A(g6488));
INVX1 NOT_340 (.Y(g7470),.A(g6927));
INVX1 NOT_341 (.Y(I15741),.A(g10260));
INVX1 NOT_342 (.Y(g7897),.A(g7712));
INVX1 NOT_343 (.Y(g7025),.A(g6400));
INVX1 NOT_344 (.Y(I6370),.A(g2356));
INVX1 NOT_345 (.Y(g7425),.A(g7214));
INVX1 NOT_346 (.Y(I11587),.A(g6828));
INVX1 NOT_347 (.Y(g2844),.A(I5966));
INVX1 NOT_348 (.Y(I12553),.A(g7676));
INVX1 NOT_349 (.Y(I12862),.A(g7638));
INVX1 NOT_350 (.Y(I8215),.A(g3981));
INVX1 NOT_351 (.Y(I10813),.A(g6397));
INVX1 NOT_352 (.Y(g11384),.A(I17209));
INVX1 NOT_353 (.Y(I14799),.A(g9661));
INVX1 NOT_354 (.Y(I6821),.A(g3015));
INVX1 NOT_355 (.Y(g2194),.A(g47));
INVX1 NOT_356 (.Y(g10160),.A(I15476));
INVX1 NOT_357 (.Y(g6797),.A(I10801));
INVX1 NOT_358 (.Y(g11067),.A(g10974));
INVX1 NOT_359 (.Y(g9342),.A(I14531));
INVX1 NOT_360 (.Y(I12326),.A(g7246));
INVX1 NOT_361 (.Y(g8928),.A(I14257));
INVX1 NOT_362 (.Y(g3121),.A(g2462));
INVX1 NOT_363 (.Y(I16280),.A(g10537));
INVX1 NOT_364 (.Y(g4160),.A(I7303));
INVX1 NOT_365 (.Y(g3321),.A(I6484));
INVX1 NOT_366 (.Y(g2089),.A(I4917));
INVX1 NOT_367 (.Y(g4933),.A(I8298));
INVX1 NOT_368 (.Y(I14973),.A(g9733));
INVX1 NOT_369 (.Y(g2731),.A(I5789));
INVX1 NOT_370 (.Y(I16688),.A(g10800));
INVX1 NOT_371 (.Y(I11543),.A(g6881));
INVX1 NOT_372 (.Y(g5420),.A(g4300));
INVX1 NOT_373 (.Y(I15801),.A(g10282));
INVX1 NOT_374 (.Y(I12948),.A(g8019));
INVX1 NOT_375 (.Y(g10455),.A(I15956));
INVX1 NOT_376 (.Y(g8064),.A(I12910));
INVX1 NOT_377 (.Y(g4521),.A(g3586));
INVX1 NOT_378 (.Y(I14805),.A(g9360));
INVX1 NOT_379 (.Y(g6291),.A(I10132));
INVX1 NOT_380 (.Y(g2557),.A(g1840));
INVX1 NOT_381 (.Y(g4050),.A(I7163));
INVX1 NOT_382 (.Y(I13117),.A(g7904));
INVX1 NOT_383 (.Y(I12904),.A(g7985));
INVX1 NOT_384 (.Y(I4873),.A(g105));
INVX1 NOT_385 (.Y(g8785),.A(I14090));
INVX1 NOT_386 (.Y(g4450),.A(g3914));
INVX1 NOT_387 (.Y(g5794),.A(I9394));
INVX1 NOT_388 (.Y(g9097),.A(g8892));
INVX1 NOT_389 (.Y(g2071),.A(I4873));
INVX1 NOT_390 (.Y(g7678),.A(I12307));
INVX1 NOT_391 (.Y(g6144),.A(I9857));
INVX1 NOT_392 (.Y(I11569),.A(g6821));
INVX1 NOT_393 (.Y(g3253),.A(I6417));
INVX1 NOT_394 (.Y(I7743),.A(g3762));
INVX1 NOT_395 (.Y(g6344),.A(I10251));
INVX1 NOT_396 (.Y(g3938),.A(g2991));
INVX1 NOT_397 (.Y(g7331),.A(I11641));
INVX1 NOT_398 (.Y(I15196),.A(g9974));
INVX1 NOT_399 (.Y(g9354),.A(I14567));
INVX1 NOT_400 (.Y(g10201),.A(g10175));
INVX1 NOT_401 (.Y(g7406),.A(I11786));
INVX1 NOT_402 (.Y(g10277),.A(I15675));
INVX1 NOT_403 (.Y(g2242),.A(I5245));
INVX1 NOT_404 (.Y(I9213),.A(g4944));
INVX1 NOT_405 (.Y(g3909),.A(g2920));
INVX1 NOT_406 (.Y(I6106),.A(g2116));
INVX1 NOT_407 (.Y(g7635),.A(I12245));
INVX1 NOT_408 (.Y(I4869),.A(g253));
INVX1 NOT_409 (.Y(I13568),.A(g8343));
INVX1 NOT_410 (.Y(I13747),.A(g8299));
INVX1 NOT_411 (.Y(I15526),.A(g10051));
INVX1 NOT_412 (.Y(g8563),.A(I13782));
INVX1 NOT_413 (.Y(g10075),.A(I15302));
INVX1 NOT_414 (.Y(g4724),.A(g3586));
INVX1 NOT_415 (.Y(g6259),.A(I10036));
INVX1 NOT_416 (.Y(g4179),.A(I7354));
INVX1 NOT_417 (.Y(g7766),.A(I12463));
INVX1 NOT_418 (.Y(I5722),.A(g2075));
INVX1 NOT_419 (.Y(g7682),.A(g7148));
INVX1 NOT_420 (.Y(I13242),.A(g8267));
INVX1 NOT_421 (.Y(I17500),.A(g11478));
INVX1 NOT_422 (.Y(g6694),.A(I10663));
INVX1 NOT_423 (.Y(g4379),.A(g3698));
INVX1 NOT_424 (.Y(g3519),.A(g3164));
INVX1 NOT_425 (.Y(g7801),.A(I12568));
INVX1 NOT_426 (.Y(g7305),.A(I11563));
INVX1 NOT_427 (.Y(I7411),.A(g4140));
INVX1 NOT_428 (.Y(g8295),.A(I13239));
INVX1 NOT_429 (.Y(g2955),.A(I6156));
INVX1 NOT_430 (.Y(I8136),.A(g4144));
INVX1 NOT_431 (.Y(g5628),.A(I9062));
INVX1 NOT_432 (.Y(I6061),.A(g2246));
INVX1 NOT_433 (.Y(I12183),.A(g7007));
INVX1 NOT_434 (.Y(g6852),.A(I10914));
INVX1 NOT_435 (.Y(I11814),.A(g7196));
INVX1 NOT_436 (.Y(g5515),.A(g4429));
INVX1 NOT_437 (.Y(I6461),.A(g2261));
INVX1 NOT_438 (.Y(g5630),.A(I9068));
INVX1 NOT_439 (.Y(I12397),.A(g7284));
INVX1 NOT_440 (.Y(I4917),.A(g584));
INVX1 NOT_441 (.Y(g2254),.A(g131));
INVX1 NOT_442 (.Y(g2814),.A(I5916));
INVX1 NOT_443 (.Y(g11402),.A(I17249));
INVX1 NOT_444 (.Y(g4289),.A(g4013));
INVX1 NOT_445 (.Y(g7748),.A(I12409));
INVX1 NOT_446 (.Y(g4777),.A(g3992));
INVX1 NOT_447 (.Y(I11807),.A(g6854));
INVX1 NOT_448 (.Y(g11457),.A(I17424));
INVX1 NOT_449 (.Y(I9090),.A(g5567));
INVX1 NOT_450 (.Y(g4835),.A(I8192));
INVX1 NOT_451 (.Y(I14400),.A(g8891));
INVX1 NOT_452 (.Y(g2350),.A(I5424));
INVX1 NOT_453 (.Y(g7755),.A(I12430));
INVX1 NOT_454 (.Y(g9267),.A(g8892));
INVX1 NOT_455 (.Y(g9312),.A(I14509));
INVX1 NOT_456 (.Y(I13639),.A(g8321));
INVX1 NOT_457 (.Y(g2038),.A(g1776));
INVX1 NOT_458 (.Y(I8943),.A(g4585));
INVX1 NOT_459 (.Y(I16763),.A(g10890));
INVX1 NOT_460 (.Y(I12933),.A(g7899));
INVX1 NOT_461 (.Y(g7226),.A(I11464));
INVX1 NOT_462 (.Y(g8089),.A(g7934));
INVX1 NOT_463 (.Y(g10352),.A(I15820));
INVX1 NOT_464 (.Y(g2438),.A(g243));
INVX1 NOT_465 (.Y(I11293),.A(g6516));
INVX1 NOT_466 (.Y(I13230),.A(g8244));
INVX1 NOT_467 (.Y(g2773),.A(I5858));
INVX1 NOT_468 (.Y(g4271),.A(g3971));
INVX1 NOT_469 (.Y(I6904),.A(g2820));
INVX1 NOT_470 (.Y(I12508),.A(g7731));
INVX1 NOT_471 (.Y(I11638),.A(g6948));
INVX1 NOT_472 (.Y(I12634),.A(g7727));
INVX1 NOT_473 (.Y(g10155),.A(I15461));
INVX1 NOT_474 (.Y(I17613),.A(g11550));
INVX1 NOT_475 (.Y(g10822),.A(I16534));
INVX1 NOT_476 (.Y(I4786),.A(g109));
INVX1 NOT_477 (.Y(I6046),.A(g2218));
INVX1 NOT_478 (.Y(I9056),.A(g4753));
INVX1 NOT_479 (.Y(g6951),.A(I11097));
INVX1 NOT_480 (.Y(g10266),.A(g10129));
INVX1 NOT_481 (.Y(I8228),.A(g4468));
INVX1 NOT_482 (.Y(I14005),.A(g8631));
INVX1 NOT_483 (.Y(g10170),.A(g10118));
INVX1 NOT_484 (.Y(I8465),.A(g4807));
INVX1 NOT_485 (.Y(I16660),.A(g10793));
INVX1 NOT_486 (.Y(g7045),.A(g6435));
INVX1 NOT_487 (.Y(I10538),.A(g5910));
INVX1 NOT_488 (.Y(I8934),.A(g4271));
INVX1 NOT_489 (.Y(I5424),.A(g910));
INVX1 NOT_490 (.Y(I5795),.A(g2462));
INVX1 NOT_491 (.Y(g7445),.A(I11845));
INVX1 NOT_492 (.Y(g6114),.A(I9795));
INVX1 NOT_493 (.Y(I5737),.A(g2100));
INVX1 NOT_494 (.Y(I6403),.A(g2337));
INVX1 NOT_495 (.Y(I5809),.A(g2356));
INVX1 NOT_496 (.Y(g6314),.A(I10201));
INVX1 NOT_497 (.Y(I7713),.A(g3750));
INVX1 NOT_498 (.Y(g9761),.A(g9454));
INVX1 NOT_499 (.Y(I11841),.A(g7226));
INVX1 NOT_500 (.Y(I11992),.A(g7058));
INVX1 NOT_501 (.Y(I11391),.A(g6387));
INVX1 NOT_502 (.Y(I9851),.A(g5405));
INVX1 NOT_503 (.Y(g2212),.A(g686));
INVX1 NOT_504 (.Y(I13391),.A(g8178));
INVX1 NOT_505 (.Y(g6870),.A(I10952));
INVX1 NOT_506 (.Y(g4674),.A(I8050));
INVX1 NOT_507 (.Y(g8948),.A(I14299));
INVX1 NOT_508 (.Y(g3141),.A(g2563));
INVX1 NOT_509 (.Y(I6391),.A(g2478));
INVX1 NOT_510 (.Y(I5672),.A(g569));
INVX1 NOT_511 (.Y(I15688),.A(g10207));
INVX1 NOT_512 (.Y(g5040),.A(I8421));
INVX1 NOT_513 (.Y(I5077),.A(g35));
INVX1 NOT_514 (.Y(g1983),.A(g750));
INVX1 NOT_515 (.Y(g6825),.A(I10873));
INVX1 NOT_516 (.Y(g3710),.A(g3215));
INVX1 NOT_517 (.Y(g7369),.A(g7273));
INVX1 NOT_518 (.Y(g7602),.A(I12156));
INVX1 NOT_519 (.Y(g10167),.A(I15497));
INVX1 NOT_520 (.Y(g10194),.A(g10062));
INVX1 NOT_521 (.Y(g10589),.A(I16252));
INVX1 NOT_522 (.Y(I16550),.A(g10726));
INVX1 NOT_523 (.Y(g4541),.A(I7946));
INVX1 NOT_524 (.Y(g7007),.A(I11146));
INVX1 NOT_525 (.Y(I17371),.A(g11410));
INVX1 NOT_526 (.Y(I17234),.A(g11353));
INVX1 NOT_527 (.Y(g7920),.A(g7516));
INVX1 NOT_528 (.Y(I11578),.A(g6824));
INVX1 NOT_529 (.Y(I12574),.A(g7522));
INVX1 NOT_530 (.Y(g10524),.A(g10458));
INVX1 NOT_531 (.Y(g2229),.A(g162));
INVX1 NOT_532 (.Y(I15157),.A(g9931));
INVX1 NOT_533 (.Y(I16307),.A(g10589));
INVX1 NOT_534 (.Y(g4332),.A(g4130));
INVX1 NOT_535 (.Y(I12205),.A(g6993));
INVX1 NOT_536 (.Y(g7767),.A(I12466));
INVX1 NOT_537 (.Y(I6159),.A(g2123));
INVX1 NOT_538 (.Y(g11157),.A(g10950));
INVX1 NOT_539 (.Y(g4680),.A(g3829));
INVX1 NOT_540 (.Y(g6136),.A(I9845));
INVX1 NOT_541 (.Y(g8150),.A(I13039));
INVX1 NOT_542 (.Y(g4209),.A(I7444));
INVX1 NOT_543 (.Y(g4353),.A(I7636));
INVX1 NOT_544 (.Y(g5666),.A(I9159));
INVX1 NOT_545 (.Y(g6336),.A(I10231));
INVX1 NOT_546 (.Y(g8350),.A(I13430));
INVX1 NOT_547 (.Y(I13586),.A(g8356));
INVX1 NOT_548 (.Y(g10119),.A(I15365));
INVX1 NOT_549 (.Y(I8337),.A(g4352));
INVX1 NOT_550 (.Y(g8438),.A(I13612));
INVX1 NOT_551 (.Y(g6594),.A(I10560));
INVX1 NOT_552 (.Y(g11066),.A(g10974));
INVX1 NOT_553 (.Y(g4802),.A(g3337));
INVX1 NOT_554 (.Y(I13442),.A(g8182));
INVX1 NOT_555 (.Y(g8009),.A(I12849));
INVX1 NOT_556 (.Y(I5304),.A(g79));
INVX1 NOT_557 (.Y(g10118),.A(I15362));
INVX1 NOT_558 (.Y(I6016),.A(g2201));
INVX1 NOT_559 (.Y(I6757),.A(g2732));
INVX1 NOT_560 (.Y(g7793),.A(I12544));
INVX1 NOT_561 (.Y(I9279),.A(g5314));
INVX1 NOT_562 (.Y(g5648),.A(I9105));
INVX1 NOT_563 (.Y(g6806),.A(I10828));
INVX1 NOT_564 (.Y(g5875),.A(g5361));
INVX1 NOT_565 (.Y(g6943),.A(I11079));
INVX1 NOT_566 (.Y(I16269),.A(g10558));
INVX1 NOT_567 (.Y(I9720),.A(g5248));
INVX1 NOT_568 (.Y(I12592),.A(g7445));
INVX1 NOT_569 (.Y(g10616),.A(I16289));
INVX1 NOT_570 (.Y(g4558),.A(g3880));
INVX1 NOT_571 (.Y(g5655),.A(I9126));
INVX1 NOT_572 (.Y(I13615),.A(g8333));
INVX1 NOT_573 (.Y(g7415),.A(I11797));
INVX1 NOT_574 (.Y(g7227),.A(I11467));
INVX1 NOT_575 (.Y(I9872),.A(g5557));
INVX1 NOT_576 (.Y(g10313),.A(I15741));
INVX1 NOT_577 (.Y(I5926),.A(g2172));
INVX1 NOT_578 (.Y(I13720),.A(g8358));
INVX1 NOT_579 (.Y(I9652),.A(g5426));
INVX1 NOT_580 (.Y(I5754),.A(g2304));
INVX1 NOT_581 (.Y(I10991),.A(g6759));
INVX1 NOT_582 (.Y(I15763),.A(g10244));
INVX1 NOT_583 (.Y(I11275),.A(g6502));
INVX1 NOT_584 (.Y(g10276),.A(I15672));
INVX1 NOT_585 (.Y(g11511),.A(I17552));
INVX1 NOT_586 (.Y(g4901),.A(I8268));
INVX1 NOT_587 (.Y(I7760),.A(g3768));
INVX1 NOT_588 (.Y(I16670),.A(g10797));
INVX1 NOT_589 (.Y(I11746),.A(g6857));
INVX1 NOT_590 (.Y(I13430),.A(g8241));
INVX1 NOT_591 (.Y(g10305),.A(I15725));
INVX1 NOT_592 (.Y(g10254),.A(g10196));
INVX1 NOT_593 (.Y(g4511),.A(g3586));
INVX1 NOT_594 (.Y(g10900),.A(I16656));
INVX1 NOT_595 (.Y(g9576),.A(I14713));
INVX1 NOT_596 (.Y(g2837),.A(g2130));
INVX1 NOT_597 (.Y(g10466),.A(I15989));
INVX1 NOT_598 (.Y(g5884),.A(I9505));
INVX1 NOT_599 (.Y(I5044),.A(g1182));
INVX1 NOT_600 (.Y(g6433),.A(I10349));
INVX1 NOT_601 (.Y(g5839),.A(I9452));
INVX1 NOT_602 (.Y(g8229),.A(g7826));
INVX1 NOT_603 (.Y(I6654),.A(g2952));
INVX1 NOT_604 (.Y(g8993),.A(I14400));
INVX1 NOT_605 (.Y(g2620),.A(g1998));
INVX1 NOT_606 (.Y(I12846),.A(g7685));
INVX1 NOT_607 (.Y(g2462),.A(I5555));
INVX1 NOT_608 (.Y(g9349),.A(I14552));
INVX1 NOT_609 (.Y(I8815),.A(g4471));
INVX1 NOT_610 (.Y(g10101),.A(I15335));
INVX1 NOT_611 (.Y(g10177),.A(I15523));
INVX1 NOT_612 (.Y(I16667),.A(g10780));
INVX1 NOT_613 (.Y(I13806),.A(g8478));
INVX1 NOT_614 (.Y(I7220),.A(g3213));
INVX1 NOT_615 (.Y(I5862),.A(g2537));
INVX1 NOT_616 (.Y(I9598),.A(g5120));
INVX1 NOT_617 (.Y(I7779),.A(g3774));
INVX1 NOT_618 (.Y(I17724),.A(g11625));
INVX1 NOT_619 (.Y(g6845),.A(I10907));
INVX1 NOT_620 (.Y(g7502),.A(I11882));
INVX1 NOT_621 (.Y(I8154),.A(g3636));
INVX1 NOT_622 (.Y(I10584),.A(g5864));
INVX1 NOT_623 (.Y(I17359),.A(g11372));
INVX1 NOT_624 (.Y(g3545),.A(I6733));
INVX1 NOT_625 (.Y(I15314),.A(g10007));
INVX1 NOT_626 (.Y(g11550),.A(I17591));
INVX1 NOT_627 (.Y(I15287),.A(g9980));
INVX1 NOT_628 (.Y(g6195),.A(g5426));
INVX1 NOT_629 (.Y(I7423),.A(g3331));
INVX1 NOT_630 (.Y(g6137),.A(I9848));
INVX1 NOT_631 (.Y(g5667),.A(I9162));
INVX1 NOT_632 (.Y(g6395),.A(I10293));
INVX1 NOT_633 (.Y(g3380),.A(I6576));
INVX1 NOT_634 (.Y(g5143),.A(g4682));
INVX1 NOT_635 (.Y(g6337),.A(I10234));
INVX1 NOT_636 (.Y(I16487),.A(g10771));
INVX1 NOT_637 (.Y(g6913),.A(I11021));
INVX1 NOT_638 (.Y(g10064),.A(I15290));
INVX1 NOT_639 (.Y(g11287),.A(g11207));
INVX1 NOT_640 (.Y(I15085),.A(g9720));
INVX1 NOT_641 (.Y(g2249),.A(g127));
INVX1 NOT_642 (.Y(I9625),.A(g5405));
INVX1 NOT_643 (.Y(g4580),.A(g3880));
INVX1 NOT_644 (.Y(I10759),.A(g5803));
INVX1 NOT_645 (.Y(g11307),.A(I17092));
INVX1 NOT_646 (.Y(g11076),.A(I16843));
INVX1 NOT_647 (.Y(I9232),.A(g4944));
INVX1 NOT_648 (.Y(g7188),.A(I11408));
INVX1 NOT_649 (.Y(g7689),.A(I12322));
INVX1 NOT_650 (.Y(I17121),.A(g11231));
INVX1 NOT_651 (.Y(g11596),.A(g11580));
INVX1 NOT_652 (.Y(g7388),.A(I11773));
INVX1 NOT_653 (.Y(I10114),.A(g5768));
INVX1 NOT_654 (.Y(I9253),.A(g5052));
INVX1 NOT_655 (.Y(I9938),.A(g5478));
INVX1 NOT_656 (.Y(g10874),.A(I16592));
INVX1 NOT_657 (.Y(g11054),.A(g10950));
INVX1 NOT_658 (.Y(g6807),.A(I10831));
INVX1 NOT_659 (.Y(I9813),.A(g5241));
INVX1 NOT_660 (.Y(I6417),.A(g2344));
INVX1 NOT_661 (.Y(g5693),.A(I9224));
INVX1 NOT_662 (.Y(g11243),.A(g11112));
INVX1 NOT_663 (.Y(I17344),.A(g11369));
INVX1 NOT_664 (.Y(g3507),.A(g3307));
INVX1 NOT_665 (.Y(g4262),.A(g4013));
INVX1 NOT_666 (.Y(g2298),.A(I5336));
INVX1 NOT_667 (.Y(g2085),.A(I4903));
INVX1 NOT_668 (.Y(I7665),.A(g3732));
INVX1 NOT_669 (.Y(g10630),.A(I16311));
INVX1 NOT_670 (.Y(g11431),.A(I17344));
INVX1 NOT_671 (.Y(g6859),.A(I10937));
INVX1 NOT_672 (.Y(g7028),.A(g6407));
INVX1 NOT_673 (.Y(I6982),.A(g2889));
INVX1 NOT_674 (.Y(g6266),.A(I10057));
INVX1 NOT_675 (.Y(I15269),.A(g9993));
INVX1 NOT_676 (.Y(g10166),.A(I15494));
INVX1 NOT_677 (.Y(g7030),.A(I11183));
INVX1 NOT_678 (.Y(I12583),.A(g7546));
INVX1 NOT_679 (.Y(I9519),.A(g4998));
INVX1 NOT_680 (.Y(g8062),.A(I12904));
INVX1 NOT_681 (.Y(g7430),.A(g7221));
INVX1 NOT_682 (.Y(I15341),.A(g10019));
INVX1 NOT_683 (.Y(I5414),.A(g904));
INVX1 NOT_684 (.Y(I16286),.A(g10540));
INVX1 NOT_685 (.Y(I7999),.A(g4114));
INVX1 NOT_686 (.Y(g2854),.A(I5986));
INVX1 NOT_687 (.Y(I17173),.A(g11293));
INVX1 NOT_688 (.Y(I5946),.A(g2176));
INVX1 NOT_689 (.Y(I10849),.A(g6734));
INVX1 NOT_690 (.Y(g11341),.A(I17146));
INVX1 NOT_691 (.Y(I7633),.A(g3474));
INVX1 NOT_692 (.Y(g4889),.A(I8240));
INVX1 NOT_693 (.Y(g2941),.A(I6118));
INVX1 NOT_694 (.Y(g6248),.A(I10003));
INVX1 NOT_695 (.Y(g11655),.A(I17767));
INVX1 NOT_696 (.Y(g9258),.A(g8892));
INVX1 NOT_697 (.Y(g3905),.A(g2920));
INVX1 NOT_698 (.Y(g10892),.A(I16638));
INVX1 NOT_699 (.Y(g9818),.A(I14955));
INVX1 NOT_700 (.Y(g9352),.A(I14561));
INVX1 NOT_701 (.Y(I7303),.A(g3262));
INVX1 NOT_702 (.Y(I8293),.A(g4779));
INVX1 NOT_703 (.Y(I10398),.A(g5820));
INVX1 NOT_704 (.Y(I13475),.A(g8173));
INVX1 NOT_705 (.Y(g11180),.A(I16941));
INVX1 NOT_706 (.Y(g7826),.A(I12627));
INVX1 NOT_707 (.Y(g3628),.A(g3111));
INVX1 NOT_708 (.Y(g6255),.A(I10024));
INVX1 NOT_709 (.Y(g4175),.A(I7342));
INVX1 NOT_710 (.Y(g6081),.A(g4977));
INVX1 NOT_711 (.Y(g6815),.A(I10855));
INVX1 NOT_712 (.Y(I10141),.A(g5683));
INVX1 NOT_713 (.Y(g4375),.A(g3638));
INVX1 NOT_714 (.Y(I10804),.A(g6388));
INVX1 NOT_715 (.Y(I5513),.A(g255));
INVX1 NOT_716 (.Y(g3630),.A(I6789));
INVX1 NOT_717 (.Y(g8788),.A(I14097));
INVX1 NOT_718 (.Y(I11222),.A(g6533));
INVX1 NOT_719 (.Y(I12282),.A(g7113));
INVX1 NOT_720 (.Y(I15335),.A(g10007));
INVX1 NOT_721 (.Y(I16601),.A(g10806));
INVX1 NOT_722 (.Y(g5113),.A(I8503));
INVX1 NOT_723 (.Y(g6692),.A(I10659));
INVX1 NOT_724 (.Y(I16187),.A(g10492));
INVX1 NOT_725 (.Y(g6097),.A(I9754));
INVX1 NOT_726 (.Y(I7732),.A(g3758));
INVX1 NOT_727 (.Y(g7910),.A(g7460));
INVX1 NOT_728 (.Y(I12357),.A(g7147));
INVX1 NOT_729 (.Y(g2219),.A(g94));
INVX1 NOT_730 (.Y(g9893),.A(I15082));
INVX1 NOT_731 (.Y(g2640),.A(g1984));
INVX1 NOT_732 (.Y(g6154),.A(I9875));
INVX1 NOT_733 (.Y(g4285),.A(g3688));
INVX1 NOT_734 (.Y(g6354),.A(g5867));
INVX1 NOT_735 (.Y(g2031),.A(g1690));
INVX1 NOT_736 (.Y(g10907),.A(I16673));
INVX1 NOT_737 (.Y(g5202),.A(g4640));
INVX1 NOT_738 (.Y(g6960),.A(I11112));
INVX1 NOT_739 (.Y(I15694),.A(g10234));
INVX1 NOT_740 (.Y(I5378),.A(g1857));
INVX1 NOT_741 (.Y(g2431),.A(I5510));
INVX1 NOT_742 (.Y(I15965),.A(g10405));
INVX1 NOT_743 (.Y(g2252),.A(I5271));
INVX1 NOT_744 (.Y(g2812),.A(g2158));
INVX1 NOT_745 (.Y(I7240),.A(g2824));
INVX1 NOT_746 (.Y(g7609),.A(I12177));
INVX1 NOT_747 (.Y(I10135),.A(g6249));
INVX1 NOT_748 (.Y(g7308),.A(I11572));
INVX1 NOT_749 (.Y(g8192),.A(I13117));
INVX1 NOT_750 (.Y(g2958),.A(I6163));
INVX1 NOT_751 (.Y(g8085),.A(g7932));
INVX1 NOT_752 (.Y(g10074),.A(I15299));
INVX1 NOT_753 (.Y(g5094),.A(I8462));
INVX1 NOT_754 (.Y(I13347),.A(g8122));
INVX1 NOT_755 (.Y(g2176),.A(g82));
INVX1 NOT_756 (.Y(g9026),.A(I14415));
INVX1 NOT_757 (.Y(g8485),.A(g8341));
INVX1 NOT_758 (.Y(g4184),.A(I7369));
INVX1 NOT_759 (.Y(g5494),.A(g4412));
INVX1 NOT_760 (.Y(g3750),.A(I6941));
INVX1 NOT_761 (.Y(g2005),.A(g928));
INVX1 NOT_762 (.Y(g7883),.A(g7689));
INVX1 NOT_763 (.Y(I7043),.A(g2908));
INVX1 NOT_764 (.Y(g4384),.A(I7707));
INVX1 NOT_765 (.Y(I9141),.A(g5402));
INVX1 NOT_766 (.Y(I9860),.A(g5405));
INVX1 NOT_767 (.Y(g5567),.A(I8982));
INVX1 NOT_768 (.Y(g4339),.A(g4144));
INVX1 NOT_769 (.Y(I9341),.A(g5013));
INVX1 NOT_770 (.Y(g10238),.A(g10191));
INVX1 NOT_771 (.Y(I16169),.A(g10448));
INVX1 NOT_772 (.Y(I9525),.A(g5001));
INVX1 NOT_773 (.Y(I14361),.A(g8951));
INVX1 NOT_774 (.Y(g2829),.A(I5943));
INVX1 NOT_775 (.Y(g11619),.A(I17675));
INVX1 NOT_776 (.Y(g2765),.A(g2184));
INVX1 NOT_777 (.Y(g9821),.A(I14964));
INVX1 NOT_778 (.Y(g11502),.A(I17525));
INVX1 NOT_779 (.Y(g7758),.A(I12439));
INVX1 NOT_780 (.Y(I5916),.A(g2217));
INVX1 NOT_781 (.Y(I13236),.A(g8245));
INVX1 NOT_782 (.Y(g7066),.A(I11275));
INVX1 NOT_783 (.Y(g7589),.A(I12099));
INVX1 NOT_784 (.Y(g4424),.A(g3688));
INVX1 NOT_785 (.Y(g3040),.A(g2135));
INVX1 NOT_786 (.Y(g4737),.A(g3440));
INVX1 NOT_787 (.Y(I11351),.A(g6698));
INVX1 NOT_788 (.Y(I13952),.A(g8451));
INVX1 NOT_789 (.Y(g5593),.A(I9013));
INVX1 NOT_790 (.Y(g6112),.A(I9789));
INVX1 NOT_791 (.Y(I13351),.A(g8214));
INVX1 NOT_792 (.Y(g6218),.A(I9965));
INVX1 NOT_793 (.Y(g6267),.A(I10060));
INVX1 NOT_794 (.Y(g3440),.A(g3041));
INVX1 NOT_795 (.Y(g6312),.A(I10195));
INVX1 NOT_796 (.Y(g11618),.A(I17672));
INVX1 NOT_797 (.Y(g9984),.A(I15184));
INVX1 NOT_798 (.Y(I11821),.A(g7205));
INVX1 NOT_799 (.Y(g10176),.A(I15520));
INVX1 NOT_800 (.Y(g10185),.A(g10040));
INVX1 NOT_801 (.Y(g10675),.A(g10574));
INVX1 NOT_802 (.Y(I16479),.A(g10767));
INVX1 NOT_803 (.Y(g10092),.A(I15323));
INVX1 NOT_804 (.Y(I10048),.A(g5734));
INVX1 NOT_805 (.Y(I16363),.A(g10599));
INVX1 NOT_806 (.Y(I16217),.A(g10501));
INVX1 NOT_807 (.Y(g3323),.A(g2157));
INVX1 NOT_808 (.Y(I15278),.A(g10033));
INVX1 NOT_809 (.Y(g7571),.A(I12035));
INVX1 NOT_810 (.Y(g7365),.A(I11743));
INVX1 NOT_811 (.Y(g2733),.A(I5795));
INVX1 NOT_812 (.Y(g4077),.A(I7202));
INVX1 NOT_813 (.Y(g6001),.A(I9625));
INVX1 NOT_814 (.Y(g7048),.A(I11225));
INVX1 NOT_815 (.Y(g10154),.A(I15458));
INVX1 NOT_816 (.Y(g2270),.A(I5311));
INVX1 NOT_817 (.Y(I5798),.A(g2085));
INVX1 NOT_818 (.Y(I17240),.A(g11395));
INVX1 NOT_819 (.Y(g7711),.A(I12344));
INVX1 NOT_820 (.Y(g4523),.A(g3546));
INVX1 NOT_821 (.Y(I10221),.A(g6117));
INVX1 NOT_822 (.Y(I11790),.A(g7246));
INVX1 NOT_823 (.Y(g8520),.A(I13729));
INVX1 NOT_824 (.Y(g6293),.A(I10138));
INVX1 NOT_825 (.Y(g11469),.A(I17444));
INVX1 NOT_826 (.Y(g8219),.A(g7826));
INVX1 NOT_827 (.Y(g2225),.A(I5210));
INVX1 NOT_828 (.Y(g8640),.A(g8512));
INVX1 NOT_829 (.Y(g10935),.A(g10827));
INVX1 NOT_830 (.Y(g2610),.A(I5731));
INVX1 NOT_831 (.Y(g2073),.A(I4879));
INVX1 NOT_832 (.Y(g2796),.A(g2276));
INVX1 NOT_833 (.Y(g11468),.A(I17441));
INVX1 NOT_834 (.Y(g11039),.A(I16778));
INVX1 NOT_835 (.Y(I6851),.A(g2937));
INVX1 NOT_836 (.Y(g4205),.A(I7432));
INVX1 NOT_837 (.Y(I7697),.A(g3743));
INVX1 NOT_838 (.Y(I10613),.A(g6000));
INVX1 NOT_839 (.Y(I11873),.A(g6863));
INVX1 NOT_840 (.Y(g10883),.A(g10809));
INVX1 NOT_841 (.Y(I17755),.A(g11646));
INVX1 NOT_842 (.Y(g7333),.A(I11647));
INVX1 NOT_843 (.Y(g9106),.A(I14439));
INVX1 NOT_844 (.Y(I7210),.A(g2798));
INVX1 NOT_845 (.Y(g7774),.A(I12487));
INVX1 NOT_846 (.Y(g5521),.A(g4530));
INVX1 NOT_847 (.Y(g3528),.A(g3164));
INVX1 NOT_848 (.Y(g8958),.A(I14323));
INVX1 NOT_849 (.Y(I16580),.A(g10826));
INVX1 NOT_850 (.Y(I17770),.A(g11649));
INVX1 NOT_851 (.Y(g11038),.A(I16775));
INVX1 NOT_852 (.Y(g5050),.A(I8429));
INVX1 NOT_853 (.Y(g2124),.A(I5050));
INVX1 NOT_854 (.Y(g3351),.A(I6535));
INVX1 NOT_855 (.Y(g5641),.A(I9084));
INVX1 NOT_856 (.Y(I17563),.A(g11492));
INVX1 NOT_857 (.Y(g2980),.A(g1983));
INVX1 NOT_858 (.Y(g6727),.A(g5997));
INVX1 NOT_859 (.Y(g8376),.A(I13478));
INVX1 NOT_860 (.Y(I5632),.A(g932));
INVX1 NOT_861 (.Y(I5095),.A(g37));
INVX1 NOT_862 (.Y(I6260),.A(g2025));
INVX1 NOT_863 (.Y(g2069),.A(I4869));
INVX1 NOT_864 (.Y(I9111),.A(g5596));
INVX1 NOT_865 (.Y(g7196),.A(I11420));
INVX1 NOT_866 (.Y(g4551),.A(g3946));
INVX1 NOT_867 (.Y(I15601),.A(g10173));
INVX1 NOT_868 (.Y(I9311),.A(g4915));
INVX1 NOT_869 (.Y(I15187),.A(g9968));
INVX1 NOT_870 (.Y(g7803),.A(I12574));
INVX1 NOT_871 (.Y(I12248),.A(g7098));
INVX1 NOT_872 (.Y(I13209),.A(g8198));
INVX1 NOT_873 (.Y(g4499),.A(g3546));
INVX1 NOT_874 (.Y(I8848),.A(g4490));
INVX1 NOT_875 (.Y(g2540),.A(I5655));
INVX1 NOT_876 (.Y(g7538),.A(I11950));
INVX1 NOT_877 (.Y(I13834),.A(g8488));
INVX1 NOT_878 (.Y(I5579),.A(g1197));
INVX1 NOT_879 (.Y(g7780),.A(I12505));
INVX1 NOT_880 (.Y(g5724),.A(I9268));
INVX1 NOT_881 (.Y(g9027),.A(I14418));
INVX1 NOT_882 (.Y(g2206),.A(I5171));
INVX1 NOT_883 (.Y(I12779),.A(g7608));
INVX1 NOT_884 (.Y(g10729),.A(g10630));
INVX1 NOT_885 (.Y(g6703),.A(I10678));
INVX1 NOT_886 (.Y(I9174),.A(g4903));
INVX1 NOT_887 (.Y(I5719),.A(g2072));
INVX1 NOT_888 (.Y(g10577),.A(g10526));
INVX1 NOT_889 (.Y(I17767),.A(g11648));
INVX1 NOT_890 (.Y(g7509),.A(I11889));
INVX1 NOT_891 (.Y(g9427),.A(g9079));
INVX1 NOT_892 (.Y(I10033),.A(g5693));
INVX1 NOT_893 (.Y(I7820),.A(g3811));
INVX1 NOT_894 (.Y(I10234),.A(g6114));
INVX1 NOT_895 (.Y(g4754),.A(g3440));
INVX1 NOT_896 (.Y(I16531),.A(g10720));
INVX1 NOT_897 (.Y(g10439),.A(g10334));
INVX1 NOT_898 (.Y(I11021),.A(g6398));
INVX1 NOT_899 (.Y(I12081),.A(g6934));
INVX1 NOT_900 (.Y(g5878),.A(g5309));
INVX1 NOT_901 (.Y(g6932),.A(I11058));
INVX1 NOT_902 (.Y(g7662),.A(I12279));
INVX1 NOT_903 (.Y(g4273),.A(g4013));
INVX1 NOT_904 (.Y(I16178),.A(g10490));
INVX1 NOT_905 (.Y(I12786),.A(g7622));
INVX1 NOT_906 (.Y(I17633),.A(g11578));
INVX1 NOT_907 (.Y(g5658),.A(I9135));
INVX1 NOT_908 (.Y(g5777),.A(I9365));
INVX1 NOT_909 (.Y(I10795),.A(g6123));
INVX1 NOT_910 (.Y(I13726),.A(g8375));
INVX1 NOT_911 (.Y(g7467),.A(g7148));
INVX1 NOT_912 (.Y(g1990),.A(g774));
INVX1 NOT_913 (.Y(I6118),.A(g2248));
INVX1 NOT_914 (.Y(g8225),.A(g7826));
INVX1 NOT_915 (.Y(I17191),.A(g11315));
INVX1 NOT_916 (.Y(I17719),.A(g11623));
INVX1 NOT_917 (.Y(I11614),.A(g6838));
INVX1 NOT_918 (.Y(g8610),.A(g8483));
INVX1 NOT_919 (.Y(I6367),.A(g2045));
INVX1 NOT_920 (.Y(I9180),.A(g4905));
INVX1 NOT_921 (.Y(I12647),.A(g7711));
INVX1 NOT_922 (.Y(I16676),.A(g10798));
INVX1 NOT_923 (.Y(I16685),.A(g10785));
INVX1 NOT_924 (.Y(I11436),.A(g6488));
INVX1 NOT_925 (.Y(I9380),.A(g5013));
INVX1 NOT_926 (.Y(g10349),.A(I15811));
INVX1 NOT_927 (.Y(g9345),.A(I14540));
INVX1 NOT_928 (.Y(I16953),.A(g11082));
INVX1 NOT_929 (.Y(I13436),.A(g8187));
INVX1 NOT_930 (.Y(I9591),.A(g5095));
INVX1 NOT_931 (.Y(I16373),.A(g10593));
INVX1 NOT_932 (.Y(g4444),.A(I7800));
INVX1 NOT_933 (.Y(g8473),.A(I13669));
INVX1 NOT_934 (.Y(g2199),.A(g48));
INVX1 NOT_935 (.Y(g11410),.A(I17271));
INVX1 NOT_936 (.Y(g2399),.A(g605));
INVX1 NOT_937 (.Y(g9763),.A(I14906));
INVX1 NOT_938 (.Y(g7093),.A(I11326));
INVX1 NOT_939 (.Y(I12999),.A(g7844));
INVX1 NOT_940 (.Y(g3372),.A(g3121));
INVX1 NOT_941 (.Y(I10514),.A(g6154));
INVX1 NOT_942 (.Y(I12380),.A(g7204));
INVX1 NOT_943 (.Y(g10906),.A(I16670));
INVX1 NOT_944 (.Y(I15479),.A(g10091));
INVX1 NOT_945 (.Y(I13320),.A(g8096));
INVX1 NOT_946 (.Y(g10083),.A(I15311));
INVX1 NOT_947 (.Y(I9020),.A(g4773));
INVX1 NOT_948 (.Y(g8124),.A(g8011));
INVX1 NOT_949 (.Y(g10284),.A(g10167));
INVX1 NOT_950 (.Y(g7256),.A(I11489));
INVX1 NOT_951 (.Y(g8980),.A(I14361));
INVX1 NOT_952 (.Y(g7816),.A(I12613));
INVX1 NOT_953 (.Y(g8324),.A(I13354));
INVX1 NOT_954 (.Y(g11479),.A(I17470));
INVX1 NOT_955 (.Y(I6193),.A(g2155));
INVX1 NOT_956 (.Y(I11593),.A(g6830));
INVX1 NOT_957 (.Y(g3143),.A(I6363));
INVX1 NOT_958 (.Y(g11363),.A(I17188));
INVX1 NOT_959 (.Y(g3343),.A(g2779));
INVX1 NOT_960 (.Y(I11122),.A(g6450));
INVX1 NOT_961 (.Y(g2797),.A(g2524));
INVX1 NOT_962 (.Y(I13122),.A(g7966));
INVX1 NOT_963 (.Y(I6549),.A(g2838));
INVX1 NOT_964 (.Y(g4543),.A(g3946));
INVX1 NOT_965 (.Y(I10421),.A(g5826));
INVX1 NOT_966 (.Y(I11464),.A(g6443));
INVX1 NOT_967 (.Y(g3566),.A(I6738));
INVX1 NOT_968 (.Y(I6971),.A(g2882));
INVX1 NOT_969 (.Y(g6716),.A(g5949));
INVX1 NOT_970 (.Y(I14421),.A(g8944));
INVX1 NOT_971 (.Y(g2245),.A(I5254));
INVX1 NOT_972 (.Y(g6149),.A(I9866));
INVX1 NOT_973 (.Y(g3988),.A(g3121));
INVX1 NOT_974 (.Y(I6686),.A(g3015));
INVX1 NOT_975 (.Y(g6349),.A(I10258));
INVX1 NOT_976 (.Y(g7847),.A(I12638));
INVX1 NOT_977 (.Y(g3693),.A(g2920));
INVX1 NOT_978 (.Y(I11034),.A(g6629));
INVX1 NOT_979 (.Y(I10012),.A(g5543));
INVX1 NOT_980 (.Y(g3334),.A(I6517));
INVX1 NOT_981 (.Y(I5725),.A(g2079));
INVX1 NOT_982 (.Y(g7685),.A(g7148));
INVX1 NOT_983 (.Y(g7197),.A(I11423));
INVX1 NOT_984 (.Y(I11641),.A(g6960));
INVX1 NOT_985 (.Y(I11797),.A(g6852));
INVX1 NOT_986 (.Y(g5997),.A(I9617));
INVX1 NOT_987 (.Y(I15580),.A(g10155));
INVX1 NOT_988 (.Y(I13797),.A(g8473));
INVX1 NOT_989 (.Y(I6598),.A(g2623));
INVX1 NOT_990 (.Y(g7021),.A(I11162));
INVX1 NOT_991 (.Y(g4729),.A(g3586));
INVX1 NOT_992 (.Y(g4961),.A(I8333));
INVX1 NOT_993 (.Y(g7421),.A(I11807));
INVX1 NOT_994 (.Y(g10139),.A(I15415));
INVX1 NOT_995 (.Y(g2344),.A(I5410));
INVX1 NOT_996 (.Y(I8211),.A(g3566));
INVX1 NOT_997 (.Y(I9905),.A(g5300));
INVX1 NOT_998 (.Y(g6398),.A(I10302));
INVX1 NOT_999 (.Y(I10541),.A(g6176));
INVX1 NOT_1000 (.Y(I6121),.A(g2121));
INVX1 NOT_1001 (.Y(g1963),.A(g110));
INVX1 NOT_1002 (.Y(I17324),.A(g11347));
INVX1 NOT_1003 (.Y(g7263),.A(I11498));
INVX1 NOT_1004 (.Y(I14473),.A(g8921));
INVX1 NOT_1005 (.Y(g2207),.A(I5174));
INVX1 NOT_1006 (.Y(g10138),.A(I15412));
INVX1 NOT_1007 (.Y(I17701),.A(g11617));
INVX1 NOT_1008 (.Y(I10789),.A(g5867));
INVX1 NOT_1009 (.Y(I12448),.A(g7530));
INVX1 NOT_1010 (.Y(I13409),.A(g8141));
INVX1 NOT_1011 (.Y(I17534),.A(g11495));
INVX1 NOT_1012 (.Y(g3792),.A(I7017));
INVX1 NOT_1013 (.Y(g5353),.A(I8820));
INVX1 NOT_1014 (.Y(g8849),.A(g8745));
INVX1 NOT_1015 (.Y(g2259),.A(I5292));
INVX1 NOT_1016 (.Y(g6241),.A(I9992));
INVX1 NOT_1017 (.Y(g2819),.A(g2159));
INVX1 NOT_1018 (.Y(I11408),.A(g6405));
INVX1 NOT_1019 (.Y(I12505),.A(g7728));
INVX1 NOT_1020 (.Y(I11635),.A(g6947));
INVX1 NOT_1021 (.Y(I10724),.A(g6096));
INVX1 NOT_1022 (.Y(g11084),.A(I16863));
INVX1 NOT_1023 (.Y(g4885),.A(I8228));
INVX1 NOT_1024 (.Y(g4414),.A(I7752));
INVX1 NOT_1025 (.Y(I10325),.A(g6003));
INVX1 NOT_1026 (.Y(g11110),.A(g10974));
INVX1 NOT_1027 (.Y(g3621),.A(I6754));
INVX1 NOT_1028 (.Y(I6938),.A(g2854));
INVX1 NOT_1029 (.Y(I7668),.A(g3733));
INVX1 NOT_1030 (.Y(g2852),.A(I5982));
INVX1 NOT_1031 (.Y(I7840),.A(g3431));
INVX1 NOT_1032 (.Y(I16543),.A(g10747));
INVX1 NOT_1033 (.Y(g10852),.A(g10740));
INVX1 NOT_1034 (.Y(g8781),.A(I14080));
INVX1 NOT_1035 (.Y(I8614),.A(g4414));
INVX1 NOT_1036 (.Y(I10920),.A(g6733));
INVX1 NOT_1037 (.Y(I10535),.A(g5867));
INVX1 NOT_1038 (.Y(I12026),.A(g7119));
INVX1 NOT_1039 (.Y(I10434),.A(g5843));
INVX1 NOT_1040 (.Y(g11179),.A(I16938));
INVX1 NOT_1041 (.Y(g2701),.A(g2040));
INVX1 NOT_1042 (.Y(g3113),.A(I6343));
INVX1 NOT_1043 (.Y(g7562),.A(g6984));
INVX1 NOT_1044 (.Y(I14358),.A(g8950));
INVX1 NOT_1045 (.Y(I7390),.A(g4087));
INVX1 NOT_1046 (.Y(I10828),.A(g6708));
INVX1 NOT_1047 (.Y(I10946),.A(g6548));
INVX1 NOT_1048 (.Y(g8797),.A(I14116));
INVX1 NOT_1049 (.Y(g6644),.A(I10601));
INVX1 NOT_1050 (.Y(g4513),.A(g3546));
INVX1 NOT_1051 (.Y(g7631),.A(I12235));
INVX1 NOT_1052 (.Y(I5171),.A(g1419));
INVX1 NOT_1053 (.Y(g7723),.A(I12354));
INVX1 NOT_1054 (.Y(g6119),.A(I9810));
INVX1 NOT_1055 (.Y(I9973),.A(g5502));
INVX1 NOT_1056 (.Y(g7817),.A(I12616));
INVX1 NOT_1057 (.Y(g5901),.A(g5361));
INVX1 NOT_1058 (.Y(I4920),.A(g260));
INVX1 NOT_1059 (.Y(g8291),.A(I13227));
INVX1 NOT_1060 (.Y(g11373),.A(I17198));
INVX1 NOT_1061 (.Y(g3094),.A(I6302));
INVX1 NOT_1062 (.Y(g6258),.A(I10033));
INVX1 NOT_1063 (.Y(g4178),.A(I7351));
INVX1 NOT_1064 (.Y(g4436),.A(g3638));
INVX1 NOT_1065 (.Y(g6818),.A(I10864));
INVX1 NOT_1066 (.Y(g4679),.A(g4013));
INVX1 NOT_1067 (.Y(g11654),.A(I17764));
INVX1 NOT_1068 (.Y(g4378),.A(I7697));
INVX1 NOT_1069 (.Y(g7605),.A(I12165));
INVX1 NOT_1070 (.Y(g5511),.A(I8934));
INVX1 NOT_1071 (.Y(I11575),.A(g6823));
INVX1 NOT_1072 (.Y(g3518),.A(g3164));
INVX1 NOT_1073 (.Y(I10682),.A(g6051));
INVX1 NOT_1074 (.Y(g10576),.A(g10524));
INVX1 NOT_1075 (.Y(I9040),.A(g4794));
INVX1 NOT_1076 (.Y(g8144),.A(I13027));
INVX1 NOT_1077 (.Y(g8344),.A(I13412));
INVX1 NOT_1078 (.Y(g6717),.A(I10706));
INVX1 NOT_1079 (.Y(I9440),.A(g5078));
INVX1 NOT_1080 (.Y(g11417),.A(I17302));
INVX1 NOT_1081 (.Y(I13711),.A(g8342));
INVX1 NOT_1082 (.Y(I16814),.A(g10910));
INVX1 NOT_1083 (.Y(I12433),.A(g7657));
INVX1 NOT_1084 (.Y(g4335),.A(I7612));
INVX1 NOT_1085 (.Y(I9123),.A(g4890));
INVX1 NOT_1086 (.Y(I11109),.A(g6464));
INVX1 NOT_1087 (.Y(g7751),.A(I12418));
INVX1 NOT_1088 (.Y(g4182),.A(I7363));
INVX1 NOT_1089 (.Y(I9323),.A(g5620));
INVX1 NOT_1090 (.Y(I13109),.A(g7981));
INVX1 NOT_1091 (.Y(g4288),.A(g4130));
INVX1 NOT_1092 (.Y(I11537),.A(g7144));
INVX1 NOT_1093 (.Y(g4382),.A(g3638));
INVX1 NOT_1094 (.Y(I16772),.A(g10887));
INVX1 NOT_1095 (.Y(g3776),.A(g2579));
INVX1 NOT_1096 (.Y(g6893),.A(I10991));
INVX1 NOT_1097 (.Y(g5574),.A(g4300));
INVX1 NOT_1098 (.Y(g5864),.A(I9483));
INVX1 NOT_1099 (.Y(g10200),.A(g10169));
INVX1 NOT_1100 (.Y(g8694),.A(I13975));
INVX1 NOT_1101 (.Y(g2825),.A(I5935));
INVX1 NOT_1102 (.Y(g2650),.A(g2006));
INVX1 NOT_1103 (.Y(g10608),.A(I16283));
INVX1 NOT_1104 (.Y(g10115),.A(I15353));
INVX1 NOT_1105 (.Y(g6386),.A(I10282));
INVX1 NOT_1106 (.Y(g7585),.A(I12081));
INVX1 NOT_1107 (.Y(I17447),.A(g11457));
INVX1 NOT_1108 (.Y(I5684),.A(g572));
INVX1 NOT_1109 (.Y(I8061),.A(g3381));
INVX1 NOT_1110 (.Y(g4805),.A(g3337));
INVX1 NOT_1111 (.Y(I7163),.A(g2643));
INVX1 NOT_1112 (.Y(I5963),.A(g2179));
INVX1 NOT_1113 (.Y(I7810),.A(g3799));
INVX1 NOT_1114 (.Y(g7041),.A(g6427));
INVX1 NOT_1115 (.Y(I7363),.A(g4005));
INVX1 NOT_1116 (.Y(I16638),.A(g10863));
INVX1 NOT_1117 (.Y(g2008),.A(g971));
INVX1 NOT_1118 (.Y(I13606),.A(g8311));
INVX1 NOT_1119 (.Y(I12971),.A(g8039));
INVX1 NOT_1120 (.Y(I11303),.A(g6526));
INVX1 NOT_1121 (.Y(g6274),.A(I10081));
INVX1 NOT_1122 (.Y(I7432),.A(g3663));
INVX1 NOT_1123 (.Y(g6426),.A(I10340));
INVX1 NOT_1124 (.Y(g11423),.A(I17324));
INVX1 NOT_1125 (.Y(g2336),.A(g1900));
INVX1 NOT_1126 (.Y(I16416),.A(g10664));
INVX1 NOT_1127 (.Y(I12369),.A(g7189));
INVX1 NOT_1128 (.Y(I9875),.A(g5278));
INVX1 NOT_1129 (.Y(I7453),.A(g3708));
INVX1 NOT_1130 (.Y(g6170),.A(g5426));
INVX1 NOT_1131 (.Y(I14506),.A(g8923));
INVX1 NOT_1132 (.Y(g7673),.A(I12296));
INVX1 NOT_1133 (.Y(I9655),.A(g5173));
INVX1 NOT_1134 (.Y(g6125),.A(I9822));
INVX1 NOT_1135 (.Y(I5707),.A(g2418));
INVX1 NOT_1136 (.Y(g8886),.A(I14228));
INVX1 NOT_1137 (.Y(g3521),.A(g3164));
INVX1 NOT_1138 (.Y(g8951),.A(I14306));
INVX1 NOT_1139 (.Y(I16510),.A(g10712));
INVX1 NOT_1140 (.Y(g5262),.A(g4353));
INVX1 NOT_1141 (.Y(g3050),.A(I6260));
INVX1 NOT_1142 (.Y(I11091),.A(g6657));
INVX1 NOT_1143 (.Y(g10973),.A(I16720));
INVX1 NOT_1144 (.Y(g5736),.A(I9296));
INVX1 NOT_1145 (.Y(g6984),.A(g6382));
INVX1 NOT_1146 (.Y(g6280),.A(I10099));
INVX1 NOT_1147 (.Y(g6939),.A(I11071));
INVX1 NOT_1148 (.Y(g7669),.A(I12286));
INVX1 NOT_1149 (.Y(I17246),.A(g11341));
INVX1 NOT_1150 (.Y(g11543),.A(g11519));
INVX1 NOT_1151 (.Y(g3996),.A(g3144));
INVX1 NOT_1152 (.Y(g10184),.A(g10039));
INVX1 NOT_1153 (.Y(I12412),.A(g7520));
INVX1 NOT_1154 (.Y(I8403),.A(g4264));
INVX1 NOT_1155 (.Y(g10674),.A(g10584));
INVX1 NOT_1156 (.Y(g8314),.A(I13326));
INVX1 NOT_1157 (.Y(g5623),.A(I9053));
INVX1 NOT_1158 (.Y(g7772),.A(I12481));
INVX1 NOT_1159 (.Y(I7157),.A(g3015));
INVX1 NOT_1160 (.Y(g7058),.A(I11255));
INVX1 NOT_1161 (.Y(I12133),.A(g6870));
INVX1 NOT_1162 (.Y(I5957),.A(g2178));
INVX1 NOT_1163 (.Y(I7357),.A(g4077));
INVX1 NOT_1164 (.Y(g2122),.A(I5044));
INVX1 NOT_1165 (.Y(g2228),.A(g28));
INVX1 NOT_1166 (.Y(g7531),.A(I11929));
INVX1 NOT_1167 (.Y(g4095),.A(I7233));
INVX1 NOT_1168 (.Y(g9554),.A(I14697));
INVX1 NOT_1169 (.Y(g8870),.A(I14182));
INVX1 NOT_1170 (.Y(g2322),.A(I5378));
INVX1 NOT_1171 (.Y(I10927),.A(g6755));
INVX1 NOT_1172 (.Y(g7458),.A(g7123));
INVX1 NOT_1173 (.Y(g5889),.A(I9514));
INVX1 NOT_1174 (.Y(I12229),.A(g7070));
INVX1 NOT_1175 (.Y(I6962),.A(g2791));
INVX1 NOT_1176 (.Y(g4495),.A(I7886));
INVX1 NOT_1177 (.Y(I9839),.A(g5226));
INVX1 NOT_1178 (.Y(g2230),.A(g704));
INVX1 NOT_1179 (.Y(g4437),.A(g3345));
INVX1 NOT_1180 (.Y(g4102),.A(I7244));
INVX1 NOT_1181 (.Y(I17591),.A(g11514));
INVX1 NOT_1182 (.Y(g4208),.A(I7441));
INVX1 NOT_1183 (.Y(g7890),.A(g7479));
INVX1 NOT_1184 (.Y(g8650),.A(I13933));
INVX1 NOT_1185 (.Y(I13840),.A(g8488));
INVX1 NOT_1186 (.Y(I16586),.A(g10850));
INVX1 NOT_1187 (.Y(g3379),.A(g3121));
INVX1 NOT_1188 (.Y(I15568),.A(g10094));
INVX1 NOT_1189 (.Y(g10934),.A(g10827));
INVX1 NOT_1190 (.Y(g6106),.A(I9773));
INVX1 NOT_1191 (.Y(g5175),.A(g4682));
INVX1 NOT_1192 (.Y(g6306),.A(I10177));
INVX1 NOT_1193 (.Y(g7505),.A(g7148));
INVX1 NOT_1194 (.Y(g3878),.A(g2920));
INVX1 NOT_1195 (.Y(g11242),.A(g11112));
INVX1 NOT_1196 (.Y(I5098),.A(g38));
INVX1 NOT_1197 (.Y(g8008),.A(I12846));
INVX1 NOT_1198 (.Y(I10240),.A(g5937));
INVX1 NOT_1199 (.Y(g7011),.A(g6503));
INVX1 NOT_1200 (.Y(g4719),.A(g3586));
INVX1 NOT_1201 (.Y(g10692),.A(I16363));
INVX1 NOT_1202 (.Y(g5651),.A(I9114));
INVX1 NOT_1203 (.Y(I6587),.A(g2620));
INVX1 NOT_1204 (.Y(I10648),.A(g6030));
INVX1 NOT_1205 (.Y(I15814),.A(g10202));
INVX1 NOT_1206 (.Y(g8336),.A(I13388));
INVX1 NOT_1207 (.Y(I14903),.A(g9507));
INVX1 NOT_1208 (.Y(I5833),.A(g2103));
INVX1 NOT_1209 (.Y(g6387),.A(g6121));
INVX1 NOT_1210 (.Y(g5285),.A(g4355));
INVX1 NOT_1211 (.Y(g6461),.A(I10391));
INVX1 NOT_1212 (.Y(I15807),.A(g10284));
INVX1 NOT_1213 (.Y(I15974),.A(g10411));
INVX1 NOT_1214 (.Y(I8858),.A(g4506));
INVX1 NOT_1215 (.Y(g2550),.A(g1834));
INVX1 NOT_1216 (.Y(g7074),.A(I11299));
INVX1 NOT_1217 (.Y(I16720),.A(g10854));
INVX1 NOT_1218 (.Y(g3271),.A(I6443));
INVX1 NOT_1219 (.Y(g10400),.A(g10348));
INVX1 NOT_1220 (.Y(g2845),.A(g2168));
INVX1 NOT_1221 (.Y(I9282),.A(g5633));
INVX1 NOT_1222 (.Y(I15639),.A(g10179));
INVX1 NOT_1223 (.Y(I10563),.A(g6043));
INVX1 NOT_1224 (.Y(I5584),.A(g1200));
INVX1 NOT_1225 (.Y(g10214),.A(I15586));
INVX1 NOT_1226 (.Y(g9490),.A(g9324));
INVX1 NOT_1227 (.Y(g9823),.A(I14970));
INVX1 NOT_1228 (.Y(g2195),.A(g83));
INVX1 NOT_1229 (.Y(g4265),.A(g3664));
INVX1 NOT_1230 (.Y(I15293),.A(g10001));
INVX1 NOT_1231 (.Y(I9988),.A(g5526));
INVX1 NOT_1232 (.Y(g6427),.A(I10343));
INVX1 NOT_1233 (.Y(I12627),.A(g7697));
INVX1 NOT_1234 (.Y(g2395),.A(g231));
INVX1 NOT_1235 (.Y(g2891),.A(I6055));
INVX1 NOT_1236 (.Y(g5184),.A(g4682));
INVX1 NOT_1237 (.Y(g2337),.A(I5395));
INVX1 NOT_1238 (.Y(I11483),.A(g6567));
INVX1 NOT_1239 (.Y(g2913),.A(I6088));
INVX1 NOT_1240 (.Y(g10329),.A(I15775));
INVX1 NOT_1241 (.Y(g10207),.A(g10186));
INVX1 NOT_1242 (.Y(g4442),.A(g3638));
INVX1 NOT_1243 (.Y(I6985),.A(g2890));
INVX1 NOT_1244 (.Y(g6904),.A(I11008));
INVX1 NOT_1245 (.Y(g6200),.A(I9935));
INVX1 NOT_1246 (.Y(g11638),.A(I17724));
INVX1 NOT_1247 (.Y(g10539),.A(I16184));
INVX1 NOT_1248 (.Y(g4786),.A(I8154));
INVX1 NOT_1249 (.Y(g6046),.A(I9669));
INVX1 NOT_1250 (.Y(g8065),.A(I12913));
INVX1 NOT_1251 (.Y(g3799),.A(I7022));
INVX1 NOT_1252 (.Y(I8315),.A(g4788));
INVX1 NOT_1253 (.Y(I8811),.A(g4465));
INVX1 NOT_1254 (.Y(g6446),.A(I10370));
INVX1 NOT_1255 (.Y(g8122),.A(I12981));
INVX1 NOT_1256 (.Y(g3981),.A(I7118));
INVX1 NOT_1257 (.Y(g8465),.A(g8289));
INVX1 NOT_1258 (.Y(g9529),.A(I14672));
INVX1 NOT_1259 (.Y(g4164),.A(I7311));
INVX1 NOT_1260 (.Y(g10538),.A(I16181));
INVX1 NOT_1261 (.Y(g4233),.A(g3698));
INVX1 NOT_1262 (.Y(g5424),.A(I8865));
INVX1 NOT_1263 (.Y(g9348),.A(I14549));
INVX1 NOT_1264 (.Y(I11326),.A(g6660));
INVX1 NOT_1265 (.Y(I13949),.A(g8451));
INVX1 NOT_1266 (.Y(g6403),.A(g6128));
INVX1 NOT_1267 (.Y(I13326),.A(g8203));
INVX1 NOT_1268 (.Y(I9804),.A(g5417));
INVX1 NOT_1269 (.Y(g6145),.A(I9860));
INVX1 NOT_1270 (.Y(g2859),.A(I5995));
INVX1 NOT_1271 (.Y(g3997),.A(I7131));
INVX1 NOT_1272 (.Y(I15510),.A(g10035));
INVX1 NOT_1273 (.Y(g9355),.A(I14570));
INVX1 NOT_1274 (.Y(I9792),.A(g5403));
INVX1 NOT_1275 (.Y(I6832),.A(g2909));
INVX1 NOT_1276 (.Y(g4454),.A(g3914));
INVX1 NOT_1277 (.Y(g8033),.A(I12875));
INVX1 NOT_1278 (.Y(g11510),.A(I17549));
INVX1 NOT_1279 (.Y(g6191),.A(g5446));
INVX1 NOT_1280 (.Y(g7569),.A(I12029));
INVX1 NOT_1281 (.Y(g5672),.A(I9177));
INVX1 NOT_1282 (.Y(g4296),.A(I7559));
INVX1 NOT_1283 (.Y(I11904),.A(g6902));
INVX1 NOT_1284 (.Y(I10633),.A(g6015));
INVX1 NOT_1285 (.Y(I10898),.A(g6735));
INVX1 NOT_1286 (.Y(g5231),.A(g4640));
INVX1 NOT_1287 (.Y(I17318),.A(g11340));
INVX1 NOT_1288 (.Y(g3332),.A(I6513));
INVX1 NOT_1289 (.Y(I11252),.A(g6542));
INVX1 NOT_1290 (.Y(g10241),.A(g10192));
INVX1 NOT_1291 (.Y(g9260),.A(g8892));
INVX1 NOT_1292 (.Y(g6695),.A(I10666));
INVX1 NOT_1293 (.Y(I10719),.A(g6003));
INVX1 NOT_1294 (.Y(I13621),.A(g8315));
INVX1 NOT_1295 (.Y(g5643),.A(I9090));
INVX1 NOT_1296 (.Y(g3353),.A(g3121));
INVX1 NOT_1297 (.Y(I7735),.A(g3759));
INVX1 NOT_1298 (.Y(I6507),.A(g2808));
INVX1 NOT_1299 (.Y(I14191),.A(g8795));
INVX1 NOT_1300 (.Y(g8096),.A(I12953));
INVX1 NOT_1301 (.Y(g2248),.A(g99));
INVX1 NOT_1302 (.Y(g11578),.A(I17616));
INVX1 NOT_1303 (.Y(g2342),.A(I5406));
INVX1 NOT_1304 (.Y(I7782),.A(g3775));
INVX1 NOT_1305 (.Y(g6107),.A(I9776));
INVX1 NOT_1306 (.Y(I17540),.A(g11498));
INVX1 NOT_1307 (.Y(I12857),.A(g7638));
INVX1 NOT_1308 (.Y(g11014),.A(I16735));
INVX1 NOT_1309 (.Y(g6307),.A(I10180));
INVX1 NOT_1310 (.Y(g3744),.A(g3307));
INVX1 NOT_1311 (.Y(g6536),.A(I10456));
INVX1 NOT_1312 (.Y(I4883),.A(g581));
INVX1 NOT_1313 (.Y(g5205),.A(g4366));
INVX1 NOT_1314 (.Y(I15586),.A(g10159));
INVX1 NOT_1315 (.Y(I8880),.A(g4537));
INVX1 NOT_1316 (.Y(g2255),.A(I5276));
INVX1 NOT_1317 (.Y(I5728),.A(g2084));
INVX1 NOT_1318 (.Y(g7688),.A(g7148));
INVX1 NOT_1319 (.Y(I12793),.A(g7619));
INVX1 NOT_1320 (.Y(g2481),.A(g882));
INVX1 NOT_1321 (.Y(I9202),.A(g4915));
INVX1 NOT_1322 (.Y(g8195),.A(I13122));
INVX1 NOT_1323 (.Y(g7976),.A(I12776));
INVX1 NOT_1324 (.Y(g8137),.A(I13010));
INVX1 NOT_1325 (.Y(g8891),.A(I14239));
INVX1 NOT_1326 (.Y(g8337),.A(I13391));
INVX1 NOT_1327 (.Y(g10235),.A(g10189));
INVX1 NOT_1328 (.Y(g4012),.A(I7154));
INVX1 NOT_1329 (.Y(I11183),.A(g6507));
INVX1 NOT_1330 (.Y(I16193),.A(g10485));
INVX1 NOT_1331 (.Y(g11442),.A(I17377));
INVX1 NOT_1332 (.Y(g2097),.A(I4935));
INVX1 NOT_1333 (.Y(I12765),.A(g7638));
INVX1 NOT_1334 (.Y(g10683),.A(g10612));
INVX1 NOT_1335 (.Y(g5742),.A(I9308));
INVX1 NOT_1336 (.Y(g2726),.A(g2021));
INVX1 NOT_1337 (.Y(g4412),.A(I7746));
INVX1 NOT_1338 (.Y(I11397),.A(g6713));
INVX1 NOT_1339 (.Y(I13397),.A(g8138));
INVX1 NOT_1340 (.Y(g2154),.A(I5067));
INVX1 NOT_1341 (.Y(g6016),.A(I9632));
INVX1 NOT_1342 (.Y(I12690),.A(g7555));
INVX1 NOT_1343 (.Y(g4189),.A(I7384));
INVX1 NOT_1344 (.Y(I5070),.A(g1194));
INVX1 NOT_1345 (.Y(g2960),.A(I6173));
INVX1 NOT_1346 (.Y(I10861),.A(g6694));
INVX1 NOT_1347 (.Y(I10573),.A(g5980));
INVX1 NOT_1348 (.Y(I9567),.A(g5556));
INVX1 NOT_1349 (.Y(g8807),.A(I14140));
INVX1 NOT_1350 (.Y(I14573),.A(g9029));
INVX1 NOT_1351 (.Y(g4888),.A(I8237));
INVX1 NOT_1352 (.Y(g7126),.A(I11367));
INVX1 NOT_1353 (.Y(I13933),.A(g8505));
INVX1 NOT_1354 (.Y(I17377),.A(g11412));
INVX1 NOT_1355 (.Y(g7326),.A(I11626));
INVX1 NOT_1356 (.Y(I10045),.A(g5727));
INVX1 NOT_1357 (.Y(g6115),.A(I9798));
INVX1 NOT_1358 (.Y(g6251),.A(I10012));
INVX1 NOT_1359 (.Y(g4171),.A(I7330));
INVX1 NOT_1360 (.Y(g6315),.A(I10204));
INVX1 NOT_1361 (.Y(g6811),.A(I10843));
INVX1 NOT_1362 (.Y(I15275),.A(g9994));
INVX1 NOT_1363 (.Y(g4371),.A(I7674));
INVX1 NOT_1364 (.Y(I14045),.A(g8603));
INVX1 NOT_1365 (.Y(I17739),.A(g11641));
INVX1 NOT_1366 (.Y(g4429),.A(I7779));
INVX1 NOT_1367 (.Y(g4787),.A(g3423));
INVX1 NOT_1368 (.Y(I8982),.A(g4728));
INVX1 NOT_1369 (.Y(g11041),.A(I16784));
INVX1 NOT_1370 (.Y(g10882),.A(I16616));
INVX1 NOT_1371 (.Y(g5754),.A(I9332));
INVX1 NOT_1372 (.Y(I9776),.A(g5353));
INVX1 NOT_1373 (.Y(I10099),.A(g5800));
INVX1 NOT_1374 (.Y(I16475),.A(g10765));
INVX1 NOT_1375 (.Y(g6447),.A(g6166));
INVX1 NOT_1376 (.Y(I10388),.A(g5830));
INVX1 NOT_1377 (.Y(I8234),.A(g4232));
INVX1 NOT_1378 (.Y(g7760),.A(I12445));
INVX1 NOT_1379 (.Y(I14388),.A(g8924));
INVX1 NOT_1380 (.Y(I8328),.A(g4801));
INVX1 NOT_1381 (.Y(I17146),.A(g11305));
INVX1 NOT_1382 (.Y(I16863),.A(g10972));
INVX1 NOT_1383 (.Y(g3092),.A(g2181));
INVX1 NOT_1384 (.Y(I14701),.A(g9291));
INVX1 NOT_1385 (.Y(I10251),.A(g6126));
INVX1 NOT_1386 (.Y(I14534),.A(g9290));
INVX1 NOT_1387 (.Y(g4281),.A(g3586));
INVX1 NOT_1388 (.Y(I9965),.A(g5493));
INVX1 NOT_1389 (.Y(g5613),.A(g4840));
INVX1 NOT_1390 (.Y(g6874),.A(I10958));
INVX1 NOT_1391 (.Y(g8142),.A(I13023));
INVX1 NOT_1392 (.Y(g2112),.A(g639));
INVX1 NOT_1393 (.Y(g8342),.A(I13406));
INVX1 NOT_1394 (.Y(g2218),.A(g85));
INVX1 NOT_1395 (.Y(I15983),.A(g10414));
INVX1 NOT_1396 (.Y(g2267),.A(I5304));
INVX1 NOT_1397 (.Y(I17698),.A(g11616));
INVX1 NOT_1398 (.Y(g11035),.A(I16766));
INVX1 NOT_1399 (.Y(g8255),.A(g7986));
INVX1 NOT_1400 (.Y(g8081),.A(g8000));
INVX1 NOT_1401 (.Y(g8481),.A(g8324));
INVX1 NOT_1402 (.Y(g2001),.A(g814));
INVX1 NOT_1403 (.Y(g7608),.A(I12174));
INVX1 NOT_1404 (.Y(g7924),.A(g7470));
INVX1 NOT_1405 (.Y(I5406),.A(g898));
INVX1 NOT_1406 (.Y(g7220),.A(I11456));
INVX1 NOT_1407 (.Y(g5572),.A(I8989));
INVX1 NOT_1408 (.Y(g5862),.A(I9479));
INVX1 NOT_1409 (.Y(I12245),.A(g7093));
INVX1 NOT_1410 (.Y(g7779),.A(I12502));
INVX1 NOT_1411 (.Y(I4780),.A(g872));
INVX1 NOT_1412 (.Y(I6040),.A(g2216));
INVX1 NOT_1413 (.Y(g6595),.A(I10563));
INVX1 NOT_1414 (.Y(g10584),.A(g10522));
INVX1 NOT_1415 (.Y(I15517),.A(g10051));
INVX1 NOT_1416 (.Y(I13574),.A(g8360));
INVX1 NOT_1417 (.Y(g2329),.A(I5383));
INVX1 NOT_1418 (.Y(g8354),.A(I13442));
INVX1 NOT_1419 (.Y(I14140),.A(g8717));
INVX1 NOT_1420 (.Y(g7023),.A(I11166));
INVX1 NOT_1421 (.Y(I7952),.A(g3664));
INVX1 NOT_1422 (.Y(g4963),.A(I8337));
INVX1 NOT_1423 (.Y(g10206),.A(g10178));
INVX1 NOT_1424 (.Y(I5801),.A(g1984));
INVX1 NOT_1425 (.Y(I7276),.A(g2861));
INVX1 NOT_1426 (.Y(g9670),.A(I14799));
INVX1 NOT_1427 (.Y(I16781),.A(g10893));
INVX1 NOT_1428 (.Y(g4791),.A(I8161));
INVX1 NOT_1429 (.Y(g7977),.A(I12779));
INVX1 NOT_1430 (.Y(g2828),.A(I5940));
INVX1 NOT_1431 (.Y(g6272),.A(I10075));
INVX1 NOT_1432 (.Y(I16236),.A(g10535));
INVX1 NOT_1433 (.Y(g3262),.A(I6432));
INVX1 NOT_1434 (.Y(g2727),.A(g2022));
INVX1 NOT_1435 (.Y(g3736),.A(I6924));
INVX1 NOT_1436 (.Y(g5534),.A(g4545));
INVX1 NOT_1437 (.Y(g5729),.A(I9279));
INVX1 NOT_1438 (.Y(g7361),.A(I11731));
INVX1 NOT_1439 (.Y(g10114),.A(I15350));
INVX1 NOT_1440 (.Y(I16175),.A(g10488));
INVX1 NOT_1441 (.Y(g9813),.A(I14948));
INVX1 NOT_1442 (.Y(I15193),.A(g9968));
INVX1 NOT_1443 (.Y(g6417),.A(g6136));
INVX1 NOT_1444 (.Y(I13051),.A(g8060));
INVX1 NOT_1445 (.Y(I15362),.A(g9987));
INVX1 NOT_1446 (.Y(g6935),.A(I11065));
INVX1 NOT_1447 (.Y(g11193),.A(g11112));
INVX1 NOT_1448 (.Y(g7051),.A(I11232));
INVX1 NOT_1449 (.Y(g10107),.A(I15341));
INVX1 NOT_1450 (.Y(I11756),.A(g7191));
INVX1 NOT_1451 (.Y(g2221),.A(I5198));
INVX1 NOT_1452 (.Y(g3076),.A(I6282));
INVX1 NOT_1453 (.Y(I13592),.A(g8362));
INVX1 NOT_1454 (.Y(g8783),.A(g8746));
INVX1 NOT_1455 (.Y(I15523),.A(g10058));
INVX1 NOT_1456 (.Y(g7327),.A(I11629));
INVX1 NOT_1457 (.Y(I12232),.A(g7072));
INVX1 NOT_1458 (.Y(I6528),.A(g3274));
INVX1 NOT_1459 (.Y(I16264),.A(g10557));
INVX1 NOT_1460 (.Y(g8979),.A(I14358));
INVX1 NOT_1461 (.Y(I16790),.A(g10900));
INVX1 NOT_1462 (.Y(I8490),.A(g4526));
INVX1 NOT_1463 (.Y(g4201),.A(I7420));
INVX1 NOT_1464 (.Y(I6648),.A(g2635));
INVX1 NOT_1465 (.Y(g8218),.A(g7826));
INVX1 NOT_1466 (.Y(I9658),.A(g5150));
INVX1 NOT_1467 (.Y(g8312),.A(I13320));
INVX1 NOT_1468 (.Y(I7546),.A(g4105));
INVX1 NOT_1469 (.Y(g6128),.A(I9829));
INVX1 NOT_1470 (.Y(g6629),.A(I10584));
INVX1 NOT_1471 (.Y(g5885),.A(g5361));
INVX1 NOT_1472 (.Y(g10345),.A(I15801));
INVX1 NOT_1473 (.Y(g7999),.A(I12825));
INVX1 NOT_1474 (.Y(g7146),.A(I11391));
INVX1 NOT_1475 (.Y(g5660),.A(I9141));
INVX1 NOT_1476 (.Y(I5445),.A(g922));
INVX1 NOT_1477 (.Y(g6330),.A(I10221));
INVX1 NOT_1478 (.Y(g7346),.A(I11686));
INVX1 NOT_1479 (.Y(I10162),.A(g5943));
INVX1 NOT_1480 (.Y(g7633),.A(I12239));
INVX1 NOT_1481 (.Y(g4049),.A(g3144));
INVX1 NOT_1482 (.Y(g3375),.A(I6569));
INVX1 NOT_1483 (.Y(g8001),.A(I12829));
INVX1 NOT_1484 (.Y(I12261),.A(g7078));
INVX1 NOT_1485 (.Y(g4449),.A(g4144));
INVX1 NOT_1486 (.Y(g3722),.A(I6894));
INVX1 NOT_1487 (.Y(I8456),.A(g4472));
INVX1 NOT_1488 (.Y(g7103),.A(I11338));
INVX1 NOT_1489 (.Y(g5903),.A(I9536));
INVX1 NOT_1490 (.Y(g4575),.A(g3880));
INVX1 NOT_1491 (.Y(g10848),.A(I16546));
INVX1 NOT_1492 (.Y(g11475),.A(I17466));
INVX1 NOT_1493 (.Y(g8293),.A(I13233));
INVX1 NOT_1494 (.Y(g8129),.A(g8015));
INVX1 NOT_1495 (.Y(I6010),.A(g2256));
INVX1 NOT_1496 (.Y(g2068),.A(I4866));
INVX1 NOT_1497 (.Y(I11152),.A(g6469));
INVX1 NOT_1498 (.Y(g8329),.A(I13367));
INVX1 NOT_1499 (.Y(g10141),.A(I15421));
INVX1 NOT_1500 (.Y(g7696),.A(g7148));
INVX1 NOT_1501 (.Y(g10804),.A(I16514));
INVX1 NOT_1502 (.Y(g6800),.A(I10810));
INVX1 NOT_1503 (.Y(g4098),.A(I7240));
INVX1 NOT_1504 (.Y(g3500),.A(I6690));
INVX1 NOT_1505 (.Y(I15437),.A(g10050));
INVX1 NOT_1506 (.Y(I16209),.A(g10452));
INVX1 NOT_1507 (.Y(I8851),.A(g4498));
INVX1 NOT_1508 (.Y(I11731),.A(g7021));
INVX1 NOT_1509 (.Y(g8828),.A(g8744));
INVX1 NOT_1510 (.Y(g11437),.A(I17362));
INVX1 NOT_1511 (.Y(g2677),.A(g2034));
INVX1 NOT_1512 (.Y(g10263),.A(g10127));
INVX1 NOT_1513 (.Y(g7753),.A(I12424));
INVX1 NOT_1514 (.Y(I9981),.A(g5514));
INVX1 NOT_1515 (.Y(g8727),.A(g8592));
INVX1 NOT_1516 (.Y(g5679),.A(I9194));
INVX1 NOT_1517 (.Y(g7508),.A(g6950));
INVX1 NOT_1518 (.Y(g3384),.A(g3143));
INVX1 NOT_1519 (.Y(g10332),.A(I15782));
INVX1 NOT_1520 (.Y(g6213),.A(g5426));
INVX1 NOT_1521 (.Y(g8592),.A(I13837));
INVX1 NOT_1522 (.Y(g7944),.A(g7410));
INVX1 NOT_1523 (.Y(I15347),.A(g9995));
INVX1 NOT_1524 (.Y(g7072),.A(I11293));
INVX1 NOT_1525 (.Y(I15253),.A(g9987));
INVX1 NOT_1526 (.Y(g10135),.A(I15403));
INVX1 NOT_1527 (.Y(I12445),.A(g7521));
INVX1 NOT_1528 (.Y(g11347),.A(I17164));
INVX1 NOT_1529 (.Y(g4896),.A(I8253));
INVX1 NOT_1530 (.Y(I7906),.A(g3907));
INVX1 NOT_1531 (.Y(g2349),.A(I5421));
INVX1 NOT_1532 (.Y(g7043),.A(I11214));
INVX1 NOT_1533 (.Y(I12499),.A(g7725));
INVX1 NOT_1534 (.Y(I11405),.A(g6627));
INVX1 NOT_1535 (.Y(g5288),.A(g4438));
INVX1 NOT_1536 (.Y(g9341),.A(I14528));
INVX1 NOT_1537 (.Y(g3424),.A(g2896));
INVX1 NOT_1538 (.Y(I9132),.A(g4893));
INVX1 NOT_1539 (.Y(g10361),.A(g10268));
INVX1 NOT_1540 (.Y(g3737),.A(g2834));
INVX1 NOT_1541 (.Y(g7443),.A(I11841));
INVX1 NOT_1542 (.Y(I9332),.A(g4935));
INVX1 NOT_1543 (.Y(g9525),.A(g9257));
INVX1 NOT_1544 (.Y(I9153),.A(g5027));
INVX1 NOT_1545 (.Y(I9680),.A(g5194));
INVX1 NOT_1546 (.Y(I10147),.A(g5697));
INVX1 NOT_1547 (.Y(I6343),.A(g1963));
INVX1 NOT_1548 (.Y(I10355),.A(g6003));
INVX1 NOT_1549 (.Y(g7116),.A(I11351));
INVX1 NOT_1550 (.Y(g5805),.A(I9409));
INVX1 NOT_1551 (.Y(g5916),.A(I9550));
INVX1 NOT_1552 (.Y(g7316),.A(I11596));
INVX1 NOT_1553 (.Y(g2198),.A(g668));
INVX1 NOT_1554 (.Y(I6282),.A(g2231));
INVX1 NOT_1555 (.Y(g4268),.A(I7523));
INVX1 NOT_1556 (.Y(I7771),.A(g3418));
INVX1 NOT_1557 (.Y(I16607),.A(g10787));
INVX1 NOT_1558 (.Y(g2855),.A(I5989));
INVX1 NOT_1559 (.Y(g4362),.A(I7651));
INVX1 NOT_1560 (.Y(I11929),.A(g6901));
INVX1 NOT_1561 (.Y(I14355),.A(g8948));
INVX1 NOT_1562 (.Y(I12989),.A(g8043));
INVX1 NOT_1563 (.Y(g11351),.A(I17170));
INVX1 NOT_1564 (.Y(g3077),.A(g2213));
INVX1 NOT_1565 (.Y(g5422),.A(g4470));
INVX1 NOT_1566 (.Y(g7034),.A(I11191));
INVX1 NOT_1567 (.Y(I10825),.A(g6588));
INVX1 NOT_1568 (.Y(g4419),.A(I7763));
INVX1 NOT_1569 (.Y(I9744),.A(g5263));
INVX1 NOT_1570 (.Y(I12056),.A(g6929));
INVX1 NOT_1571 (.Y(I10370),.A(g5857));
INVX1 NOT_1572 (.Y(g6166),.A(I9893));
INVX1 NOT_1573 (.Y(g8624),.A(g8486));
INVX1 NOT_1574 (.Y(g3523),.A(g2971));
INVX1 NOT_1575 (.Y(I14370),.A(g8954));
INVX1 NOT_1576 (.Y(g8953),.A(I14312));
INVX1 NOT_1577 (.Y(I10858),.A(g6688));
INVX1 NOT_1578 (.Y(I13020),.A(g8049));
INVX1 NOT_1579 (.Y(I13583),.A(g8344));
INVX1 NOT_1580 (.Y(g4452),.A(g3365));
INVX1 NOT_1581 (.Y(I8872),.A(g4529));
INVX1 NOT_1582 (.Y(I15063),.A(g9699));
INVX1 NOT_1583 (.Y(g2241),.A(g722));
INVX1 NOT_1584 (.Y(g7147),.A(I11394));
INVX1 NOT_1585 (.Y(g6056),.A(g5426));
INVX1 NOT_1586 (.Y(g5947),.A(I9585));
INVX1 NOT_1587 (.Y(g7347),.A(I11689));
INVX1 NOT_1588 (.Y(g11063),.A(g10974));
INVX1 NOT_1589 (.Y(I11046),.A(g6635));
INVX1 NOT_1590 (.Y(I10996),.A(g6786));
INVX1 NOT_1591 (.Y(I12271),.A(g7218));
INVX1 NOT_1592 (.Y(g7681),.A(g7148));
INVX1 NOT_1593 (.Y(g6649),.A(I10610));
INVX1 NOT_1594 (.Y(I8989),.A(g4746));
INVX1 NOT_1595 (.Y(g8677),.A(I13962));
INVX1 NOT_1596 (.Y(g110),.A(I4786));
INVX1 NOT_1597 (.Y(I10367),.A(g6234));
INVX1 NOT_1598 (.Y(I10394),.A(g5824));
INVX1 NOT_1599 (.Y(I9901),.A(g5557));
INVX1 NOT_1600 (.Y(g7697),.A(g7101));
INVX1 NOT_1601 (.Y(I14367),.A(g8953));
INVX1 NOT_1602 (.Y(I14394),.A(g8884));
INVX1 NOT_1603 (.Y(I16641),.A(g10864));
INVX1 NOT_1604 (.Y(g3742),.A(I6929));
INVX1 NOT_1605 (.Y(g7914),.A(g7651));
INVX1 NOT_1606 (.Y(g8576),.A(I13819));
INVX1 NOT_1607 (.Y(g2524),.A(g986));
INVX1 NOT_1608 (.Y(g7210),.A(I11440));
INVX1 NOT_1609 (.Y(g4728),.A(I8080));
INVX1 NOT_1610 (.Y(I16292),.A(g10551));
INVX1 NOT_1611 (.Y(g2644),.A(g1990));
INVX1 NOT_1612 (.Y(g6698),.A(I10671));
INVX1 NOT_1613 (.Y(g4730),.A(g3546));
INVX1 NOT_1614 (.Y(g8716),.A(g8576));
INVX1 NOT_1615 (.Y(I17546),.A(g11500));
INVX1 NOT_1616 (.Y(g8149),.A(I13036));
INVX1 NOT_1617 (.Y(g10947),.A(I16708));
INVX1 NOT_1618 (.Y(g4504),.A(I7899));
INVX1 NOT_1619 (.Y(I11357),.A(g6594));
INVX1 NOT_1620 (.Y(g6964),.A(g6509));
INVX1 NOT_1621 (.Y(g8349),.A(I13427));
INVX1 NOT_1622 (.Y(g2119),.A(I5031));
INVX1 NOT_1623 (.Y(g5095),.A(I8465));
INVX1 NOT_1624 (.Y(g6260),.A(I10039));
INVX1 NOT_1625 (.Y(g5037),.A(I8414));
INVX1 NOT_1626 (.Y(I13357),.A(g8125));
INVX1 NOT_1627 (.Y(I12199),.A(g7278));
INVX1 NOT_1628 (.Y(g4185),.A(I7372));
INVX1 NOT_1629 (.Y(I7244),.A(g3226));
INVX1 NOT_1630 (.Y(g9311),.A(I14506));
INVX1 NOT_1631 (.Y(g11422),.A(I17321));
INVX1 NOT_1632 (.Y(I11743),.A(g7035));
INVX1 NOT_1633 (.Y(I13105),.A(g7929));
INVX1 NOT_1634 (.Y(g5653),.A(I9120));
INVX1 NOT_1635 (.Y(g4385),.A(I7710));
INVX1 NOT_1636 (.Y(g7413),.A(g7197));
INVX1 NOT_1637 (.Y(g5102),.A(I8476));
INVX1 NOT_1638 (.Y(g2258),.A(I5289));
INVX1 NOT_1639 (.Y(I14319),.A(g8816));
INVX1 NOT_1640 (.Y(g2352),.A(I5430));
INVX1 NOT_1641 (.Y(g2818),.A(I5922));
INVX1 NOT_1642 (.Y(I7140),.A(g2641));
INVX1 NOT_1643 (.Y(g6063),.A(g5446));
INVX1 NOT_1644 (.Y(I12529),.A(g7589));
INVX1 NOT_1645 (.Y(I5940),.A(g2175));
INVX1 NOT_1646 (.Y(g2867),.A(I6007));
INVX1 NOT_1647 (.Y(I16635),.A(g10862));
INVX1 NOT_1648 (.Y(g10463),.A(I15980));
INVX1 NOT_1649 (.Y(g11208),.A(g11077));
INVX1 NOT_1650 (.Y(g4470),.A(I7843));
INVX1 NOT_1651 (.Y(g8198),.A(I13131));
INVX1 NOT_1652 (.Y(g4897),.A(I8256));
INVX1 NOT_1653 (.Y(g8747),.A(I14040));
INVX1 NOT_1654 (.Y(I7478),.A(g3566));
INVX1 NOT_1655 (.Y(g5719),.A(I9259));
INVX1 NOT_1656 (.Y(g4425),.A(I7771));
INVX1 NOT_1657 (.Y(I12843),.A(g7683));
INVX1 NOT_1658 (.Y(I15542),.A(g10065));
INVX1 NOT_1659 (.Y(g10972),.A(I16717));
INVX1 NOT_1660 (.Y(g10033),.A(I15235));
INVX1 NOT_1661 (.Y(I5388),.A(g889));
INVX1 NOT_1662 (.Y(g10234),.A(g10188));
INVX1 NOT_1663 (.Y(I7435),.A(g3459));
INVX1 NOT_1664 (.Y(g7936),.A(g7712));
INVX1 NOT_1665 (.Y(g11542),.A(g11519));
INVX1 NOT_1666 (.Y(g11453),.A(I17416));
INVX1 NOT_1667 (.Y(g5752),.A(I9326));
INVX1 NOT_1668 (.Y(I6094),.A(g2110));
INVX1 NOT_1669 (.Y(I13803),.A(g8476));
INVX1 NOT_1670 (.Y(g3044),.A(I6256));
INVX1 NOT_1671 (.Y(g2211),.A(g153));
INVX1 NOT_1672 (.Y(I14540),.A(g9310));
INVX1 NOT_1673 (.Y(g6279),.A(I10096));
INVX1 NOT_1674 (.Y(g2186),.A(g90));
INVX1 NOT_1675 (.Y(g7317),.A(I11599));
INVX1 NOT_1676 (.Y(g6720),.A(I10713));
INVX1 NOT_1677 (.Y(I8253),.A(g4637));
INVX1 NOT_1678 (.Y(g6118),.A(I9807));
INVX1 NOT_1679 (.Y(g3983),.A(g3222));
INVX1 NOT_1680 (.Y(g11614),.A(I17662));
INVX1 NOT_1681 (.Y(g7601),.A(I12153));
INVX1 NOT_1682 (.Y(I5430),.A(g916));
INVX1 NOT_1683 (.Y(g5265),.A(g4362));
INVX1 NOT_1684 (.Y(g11436),.A(I17359));
INVX1 NOT_1685 (.Y(g3862),.A(g2920));
INVX1 NOT_1686 (.Y(g5042),.A(g4840));
INVX1 NOT_1687 (.Y(I15320),.A(g10013));
INVX1 NOT_1688 (.Y(g9832),.A(I14989));
INVX1 NOT_1689 (.Y(g6652),.A(I10613));
INVX1 NOT_1690 (.Y(g4678),.A(g3546));
INVX1 NOT_1691 (.Y(g6057),.A(g5446));
INVX1 NOT_1692 (.Y(g6843),.A(I10901));
INVX1 NOT_1693 (.Y(I15530),.A(g10107));
INVX1 NOT_1694 (.Y(g11073),.A(g10913));
INVX1 NOT_1695 (.Y(g4331),.A(I7606));
INVX1 NOT_1696 (.Y(g3543),.A(g3101));
INVX1 NOT_1697 (.Y(g2170),.A(g30));
INVX1 NOT_1698 (.Y(g2614),.A(g1994));
INVX1 NOT_1699 (.Y(g7775),.A(I12490));
INVX1 NOT_1700 (.Y(g11593),.A(I17633));
INVX1 NOT_1701 (.Y(g7922),.A(I12712));
INVX1 NOT_1702 (.Y(g2125),.A(I5053));
INVX1 NOT_1703 (.Y(g8319),.A(I13341));
INVX1 NOT_1704 (.Y(g11346),.A(I17161));
INVX1 NOT_1705 (.Y(I15565),.A(g10101));
INVX1 NOT_1706 (.Y(g2821),.A(I5929));
INVX1 NOT_1707 (.Y(g9507),.A(g9268));
INVX1 NOT_1708 (.Y(I15464),.A(g10094));
INVX1 NOT_1709 (.Y(I6965),.A(g2880));
INVX1 NOT_1710 (.Y(I10120),.A(g6248));
INVX1 NOT_1711 (.Y(g4766),.A(g3440));
INVX1 NOT_1712 (.Y(I11662),.A(g7033));
INVX1 NOT_1713 (.Y(I10739),.A(g5942));
INVX1 NOT_1714 (.Y(g4087),.A(I7220));
INVX1 NOT_1715 (.Y(g4105),.A(I7249));
INVX1 NOT_1716 (.Y(g8152),.A(I13043));
INVX1 NOT_1717 (.Y(g10421),.A(g10331));
INVX1 NOT_1718 (.Y(I16537),.A(g10721));
INVX1 NOT_1719 (.Y(g8352),.A(I13436));
INVX1 NOT_1720 (.Y(g4305),.A(g4013));
INVX1 NOT_1721 (.Y(g6971),.A(g6517));
INVX1 NOT_1722 (.Y(I13027),.A(g8051));
INVX1 NOT_1723 (.Y(I12258),.A(g7103));
INVX1 NOT_1724 (.Y(g3729),.A(I6907));
INVX1 NOT_1725 (.Y(I6264),.A(g2118));
INVX1 NOT_1726 (.Y(I16108),.A(g10383));
INVX1 NOT_1727 (.Y(g6686),.A(I10651));
INVX1 NOT_1728 (.Y(g10163),.A(I15485));
INVX1 NOT_1729 (.Y(g8717),.A(I14010));
INVX1 NOT_1730 (.Y(g11034),.A(I16763));
INVX1 NOT_1731 (.Y(g7460),.A(g7148));
INVX1 NOT_1732 (.Y(g7597),.A(I12133));
INVX1 NOT_1733 (.Y(g5296),.A(g4444));
INVX1 NOT_1734 (.Y(I11249),.A(g6541));
INVX1 NOT_1735 (.Y(I5638),.A(g936));
INVX1 NOT_1736 (.Y(I14645),.A(g9088));
INVX1 NOT_1737 (.Y(I16283),.A(g10538));
INVX1 NOT_1738 (.Y(g2083),.A(g139));
INVX1 NOT_1739 (.Y(I6360),.A(g2261));
INVX1 NOT_1740 (.Y(g4748),.A(g3546));
INVX1 NOT_1741 (.Y(I16492),.A(g10773));
INVX1 NOT_1742 (.Y(I13482),.A(g8193));
INVX1 NOT_1743 (.Y(I5308),.A(g97));
INVX1 NOT_1744 (.Y(I11710),.A(g7020));
INVX1 NOT_1745 (.Y(g7784),.A(I12517));
INVX1 NOT_1746 (.Y(I4992),.A(g1170));
INVX1 NOT_1747 (.Y(g4755),.A(g3440));
INVX1 NOT_1748 (.Y(g10541),.A(I16190));
INVX1 NOT_1749 (.Y(I10698),.A(g5856));
INVX1 NOT_1750 (.Y(g6121),.A(I9816));
INVX1 NOT_1751 (.Y(I15409),.A(g10065));
INVX1 NOT_1752 (.Y(I7002),.A(g2907));
INVX1 NOT_1753 (.Y(g8186),.A(I13109));
INVX1 NOT_1754 (.Y(g10473),.A(g10380));
INVX1 NOT_1755 (.Y(g4226),.A(g3698));
INVX1 NOT_1756 (.Y(I11204),.A(g6523));
INVX1 NOT_1757 (.Y(g6670),.A(I10633));
INVX1 NOT_1758 (.Y(I7402),.A(g4121));
INVX1 NOT_1759 (.Y(g11409),.A(I17268));
INVX1 NOT_1760 (.Y(I6996),.A(g2904));
INVX1 NOT_1761 (.Y(g3946),.A(I7099));
INVX1 NOT_1762 (.Y(I13779),.A(g8514));
INVX1 NOT_1763 (.Y(I7236),.A(g3219));
INVX1 NOT_1764 (.Y(I15635),.A(g10185));
INVX1 NOT_1765 (.Y(I16982),.A(g11088));
INVX1 NOT_1766 (.Y(g8599),.A(g8546));
INVX1 NOT_1767 (.Y(g7995),.A(I12817));
INVX1 NOT_1768 (.Y(g2790),.A(g2276));
INVX1 NOT_1769 (.Y(g11408),.A(I17265));
INVX1 NOT_1770 (.Y(g7079),.A(I11312));
INVX1 NOT_1771 (.Y(g11635),.A(I17719));
INVX1 NOT_1772 (.Y(I11778),.A(g7210));
INVX1 NOT_1773 (.Y(g3903),.A(I7070));
INVX1 NOT_1774 (.Y(g5012),.A(I8388));
INVX1 NOT_1775 (.Y(g9100),.A(g8892));
INVX1 NOT_1776 (.Y(g8274),.A(I13194));
INVX1 NOT_1777 (.Y(I10427),.A(g5839));
INVX1 NOT_1778 (.Y(g7479),.A(I11873));
INVX1 NOT_1779 (.Y(g8426),.A(I13592));
INVX1 NOT_1780 (.Y(g1994),.A(g794));
INVX1 NOT_1781 (.Y(g4445),.A(I7803));
INVX1 NOT_1782 (.Y(g6253),.A(I10018));
INVX1 NOT_1783 (.Y(g2061),.A(g1828));
INVX1 NOT_1784 (.Y(g2187),.A(g746));
INVX1 NOT_1785 (.Y(g6938),.A(I11068));
INVX1 NOT_1786 (.Y(g4173),.A(I7336));
INVX1 NOT_1787 (.Y(g6813),.A(I10849));
INVX1 NOT_1788 (.Y(g4373),.A(I7680));
INVX1 NOT_1789 (.Y(I11786),.A(g7246));
INVX1 NOT_1790 (.Y(I16796),.A(g11016));
INVX1 NOT_1791 (.Y(g10535),.A(I16172));
INVX1 NOT_1792 (.Y(g4491),.A(g3546));
INVX1 NOT_1793 (.Y(g8125),.A(I12986));
INVX1 NOT_1794 (.Y(g7190),.A(I11412));
INVX1 NOT_1795 (.Y(g8325),.A(I13357));
INVX1 NOT_1796 (.Y(I11647),.A(g6925));
INVX1 NOT_1797 (.Y(g7390),.A(g6847));
INVX1 NOT_1798 (.Y(I12878),.A(g7638));
INVX1 NOT_1799 (.Y(g5888),.A(g5102));
INVX1 NOT_1800 (.Y(I13945),.A(g8488));
INVX1 NOT_1801 (.Y(I12171),.A(g6885));
INVX1 NOT_1802 (.Y(g10121),.A(I15371));
INVX1 NOT_1803 (.Y(g8984),.A(I14373));
INVX1 NOT_1804 (.Y(g3436),.A(g3144));
INVX1 NOT_1805 (.Y(g4369),.A(I7668));
INVX1 NOT_1806 (.Y(g8280),.A(I13212));
INVX1 NOT_1807 (.Y(I7556),.A(g4080));
INVX1 NOT_1808 (.Y(g4602),.A(I8011));
INVX1 NOT_1809 (.Y(g7501),.A(I11879));
INVX1 NOT_1810 (.Y(I17450),.A(g11450));
INVX1 NOT_1811 (.Y(g3378),.A(I6572));
INVX1 NOT_1812 (.Y(g5787),.A(I9383));
INVX1 NOT_1813 (.Y(I9424),.A(g4963));
INVX1 NOT_1814 (.Y(I9795),.A(g5404));
INVX1 NOT_1815 (.Y(I17315),.A(g11393));
INVX1 NOT_1816 (.Y(g10344),.A(I15798));
INVX1 NOT_1817 (.Y(I9737),.A(g5258));
INVX1 NOT_1818 (.Y(g2904),.A(I6065));
INVX1 NOT_1819 (.Y(g2200),.A(g92));
INVX1 NOT_1820 (.Y(g6552),.A(g5733));
INVX1 NOT_1821 (.Y(g7356),.A(I11716));
INVX1 NOT_1822 (.Y(g2046),.A(g1845));
INVX1 NOT_1823 (.Y(I17707),.A(g11619));
INVX1 NOT_1824 (.Y(g4920),.A(I8293));
INVX1 NOT_1825 (.Y(I5827),.A(g2271));
INVX1 NOT_1826 (.Y(g2446),.A(g1400));
INVX1 NOT_1827 (.Y(g4459),.A(I7820));
INVX1 NOT_1828 (.Y(I17202),.A(g11322));
INVX1 NOT_1829 (.Y(g3335),.A(I6520));
INVX1 NOT_1830 (.Y(I13233),.A(g8265));
INVX1 NOT_1831 (.Y(g8483),.A(g8332));
INVX1 NOT_1832 (.Y(g4767),.A(I8123));
INVX1 NOT_1833 (.Y(I7064),.A(g2984));
INVX1 NOT_1834 (.Y(g11575),.A(g11561));
INVX1 NOT_1835 (.Y(g2003),.A(g822));
INVX1 NOT_1836 (.Y(g5281),.A(g4428));
INVX1 NOT_1837 (.Y(g3382),.A(I6580));
INVX1 NOT_1838 (.Y(I9077),.A(g4765));
INVX1 NOT_1839 (.Y(I7899),.A(g3380));
INVX1 NOT_1840 (.Y(g4535),.A(g3946));
INVX1 NOT_1841 (.Y(I8358),.A(g4794));
INVX1 NOT_1842 (.Y(I6611),.A(g2626));
INVX1 NOT_1843 (.Y(I8506),.A(g4334));
INVX1 NOT_1844 (.Y(g2345),.A(g1936));
INVX1 NOT_1845 (.Y(g10173),.A(g10120));
INVX1 NOT_1846 (.Y(I17070),.A(g11233));
INVX1 NOT_1847 (.Y(g8106),.A(g7950));
INVX1 NOT_1848 (.Y(g11109),.A(g10974));
INVX1 NOT_1849 (.Y(g8306),.A(I13290));
INVX1 NOT_1850 (.Y(g2763),.A(I5847));
INVX1 NOT_1851 (.Y(g2191),.A(g1696));
INVX1 NOT_1852 (.Y(g2391),.A(I5478));
INVX1 NOT_1853 (.Y(g6586),.A(g5949));
INVX1 NOT_1854 (.Y(I12919),.A(g8003));
INVX1 NOT_1855 (.Y(I6799),.A(g2750));
INVX1 NOT_1856 (.Y(I11932),.A(g6908));
INVX1 NOT_1857 (.Y(g3749),.A(I6938));
INVX1 NOT_1858 (.Y(g8790),.A(I14101));
INVX1 NOT_1859 (.Y(I9205),.A(g5309));
INVX1 NOT_1860 (.Y(g11108),.A(g10974));
INVX1 NOT_1861 (.Y(g2695),.A(g2039));
INVX1 NOT_1862 (.Y(g9666),.A(I14793));
INVX1 NOT_1863 (.Y(g8061),.A(I12901));
INVX1 NOT_1864 (.Y(g5684),.A(I9205));
INVX1 NOT_1865 (.Y(I8275),.A(g4351));
INVX1 NOT_1866 (.Y(I8311),.A(g4794));
INVX1 NOT_1867 (.Y(g4415),.A(g3914));
INVX1 NOT_1868 (.Y(g5639),.A(I9080));
INVX1 NOT_1869 (.Y(I14127),.A(g8768));
INVX1 NOT_1870 (.Y(I17384),.A(g11437));
INVX1 NOT_1871 (.Y(g7810),.A(I12595));
INVX1 NOT_1872 (.Y(g7363),.A(I11737));
INVX1 NOT_1873 (.Y(g10134),.A(I15400));
INVX1 NOT_1874 (.Y(I7295),.A(g3260));
INVX1 NOT_1875 (.Y(I11961),.A(g7053));
INVX1 NOT_1876 (.Y(I16553),.A(g10754));
INVX1 NOT_1877 (.Y(g5109),.A(I8495));
INVX1 NOT_1878 (.Y(g5791),.A(I9391));
INVX1 NOT_1879 (.Y(g3798),.A(g3228));
INVX1 NOT_1880 (.Y(I13448),.A(g8150));
INVX1 NOT_1881 (.Y(I9099),.A(g5572));
INVX1 NOT_1882 (.Y(g2159),.A(I5080));
INVX1 NOT_1883 (.Y(g7432),.A(I11824));
INVX1 NOT_1884 (.Y(I14490),.A(g8885));
INVX1 NOT_1885 (.Y(g6141),.A(I9854));
INVX1 NOT_1886 (.Y(g8622),.A(g8485));
INVX1 NOT_1887 (.Y(g6570),.A(g5949));
INVX1 NOT_1888 (.Y(g6860),.A(g6475));
INVX1 NOT_1889 (.Y(g7053),.A(I11238));
INVX1 NOT_1890 (.Y(I11505),.A(g6585));
INVX1 NOT_1891 (.Y(g9351),.A(I14558));
INVX1 NOT_1892 (.Y(I5662),.A(g563));
INVX1 NOT_1893 (.Y(g9875),.A(I15036));
INVX1 NOT_1894 (.Y(g8427),.A(I13595));
INVX1 NOT_1895 (.Y(I5067),.A(g33));
INVX1 NOT_1896 (.Y(g9530),.A(I14675));
INVX1 NOT_1897 (.Y(g6710),.A(I10693));
INVX1 NOT_1898 (.Y(g5808),.A(g5320));
INVX1 NOT_1899 (.Y(I5418),.A(g907));
INVX1 NOT_1900 (.Y(g2858),.A(I5992));
INVX1 NOT_1901 (.Y(I12598),.A(g7628));
INVX1 NOT_1902 (.Y(I7194),.A(g2629));
INVX1 NOT_1903 (.Y(I14376),.A(g8959));
INVX1 NOT_1904 (.Y(I14385),.A(g8890));
INVX1 NOT_1905 (.Y(g4203),.A(I7426));
INVX1 NOT_1906 (.Y(I8985),.A(g4733));
INVX1 NOT_1907 (.Y(I13717),.A(g8354));
INVX1 NOT_1908 (.Y(g11381),.A(I17206));
INVX1 NOT_1909 (.Y(g4721),.A(g3546));
INVX1 NOT_1910 (.Y(g2016),.A(g1361));
INVX1 NOT_1911 (.Y(I13212),.A(g8195));
INVX1 NOT_1912 (.Y(g2757),.A(I5837));
INVX1 NOT_1913 (.Y(g8446),.A(I13636));
INVX1 NOT_1914 (.Y(g7568),.A(I12026));
INVX1 NOT_1915 (.Y(g5759),.A(I9341));
INVX1 NOT_1916 (.Y(I9754),.A(g5271));
INVX1 NOT_1917 (.Y(I10888),.A(g6333));
INVX1 NOT_1918 (.Y(g8514),.A(I13711));
INVX1 NOT_1919 (.Y(I6802),.A(g2751));
INVX1 NOT_1920 (.Y(g3632),.A(I6799));
INVX1 NOT_1921 (.Y(g3095),.A(g2482));
INVX1 NOT_1922 (.Y(g3037),.A(g2135));
INVX1 NOT_1923 (.Y(g8003),.A(I12835));
INVX1 NOT_1924 (.Y(I14888),.A(g9454));
INVX1 NOT_1925 (.Y(I16252),.A(g10515));
INVX1 NOT_1926 (.Y(g3437),.A(I6654));
INVX1 NOT_1927 (.Y(I12817),.A(g7692));
INVX1 NOT_1928 (.Y(I9273),.A(g5091));
INVX1 NOT_1929 (.Y(I10671),.A(g6045));
INVX1 NOT_1930 (.Y(I17695),.A(g11614));
INVX1 NOT_1931 (.Y(g3102),.A(g2482));
INVX1 NOT_1932 (.Y(I4924),.A(g123));
INVX1 NOT_1933 (.Y(g3208),.A(I6381));
INVX1 NOT_1934 (.Y(I12322),.A(g7246));
INVX1 NOT_1935 (.Y(g7912),.A(g7651));
INVX1 NOT_1936 (.Y(g8145),.A(I13030));
INVX1 NOT_1937 (.Y(g8345),.A(I13415));
INVX1 NOT_1938 (.Y(g2251),.A(g731));
INVX1 NOT_1939 (.Y(g2642),.A(g1988));
INVX1 NOT_1940 (.Y(I12159),.A(g7243));
INVX1 NOT_1941 (.Y(g7357),.A(I11719));
INVX1 NOT_1942 (.Y(g2047),.A(g1857));
INVX1 NOT_1943 (.Y(I12532),.A(g7594));
INVX1 NOT_1944 (.Y(I12901),.A(g7984));
INVX1 NOT_1945 (.Y(g8191),.A(I13114));
INVX1 NOT_1946 (.Y(g10927),.A(g10827));
INVX1 NOT_1947 (.Y(g9884),.A(I15063));
INVX1 NOT_1948 (.Y(g6158),.A(I9883));
INVX1 NOT_1949 (.Y(g3719),.A(g2920));
INVX1 NOT_1950 (.Y(I12783),.A(g7590));
INVX1 NOT_1951 (.Y(g11390),.A(I17219));
INVX1 NOT_1952 (.Y(I13723),.A(g8359));
INVX1 NOT_1953 (.Y(g5865),.A(I9486));
INVX1 NOT_1954 (.Y(g8695),.A(I13978));
INVX1 NOT_1955 (.Y(I5847),.A(g2275));
INVX1 NOT_1956 (.Y(I6901),.A(g2818));
INVX1 NOT_1957 (.Y(I11149),.A(g6468));
INVX1 NOT_1958 (.Y(g2874),.A(I6022));
INVX1 NOT_1959 (.Y(g7929),.A(g7519));
INVX1 NOT_1960 (.Y(g3752),.A(I6947));
INVX1 NOT_1961 (.Y(I16673),.A(g10782));
INVX1 NOT_1962 (.Y(I11433),.A(g6424));
INVX1 NOT_1963 (.Y(I16847),.A(g10886));
INVX1 NOT_1964 (.Y(I11387),.A(g6672));
INVX1 NOT_1965 (.Y(g5604),.A(I9032));
INVX1 NOT_1966 (.Y(I13433),.A(g8181));
INVX1 NOT_1967 (.Y(g5098),.A(g4840));
INVX1 NOT_1968 (.Y(g2654),.A(g2012));
INVX1 NOT_1969 (.Y(I11620),.A(g6840));
INVX1 NOT_1970 (.Y(g4188),.A(I7381));
INVX1 NOT_1971 (.Y(g5498),.A(I8919));
INVX1 NOT_1972 (.Y(I9712),.A(g5230));
INVX1 NOT_1973 (.Y(g6587),.A(g5827));
INVX1 NOT_1974 (.Y(g4388),.A(I7719));
INVX1 NOT_1975 (.Y(g10491),.A(I16108));
INVX1 NOT_1976 (.Y(g10903),.A(g10809));
INVX1 NOT_1977 (.Y(I11097),.A(g6748));
INVX1 NOT_1978 (.Y(I5421),.A(g549));
INVX1 NOT_1979 (.Y(g8359),.A(I13457));
INVX1 NOT_1980 (.Y(g6111),.A(I9786));
INVX1 NOT_1981 (.Y(g6275),.A(I10084));
INVX1 NOT_1982 (.Y(g6311),.A(I10192));
INVX1 NOT_1983 (.Y(g4216),.A(I7465));
INVX1 NOT_1984 (.Y(g10604),.A(I16280));
INVX1 NOT_1985 (.Y(g9343),.A(I14534));
INVX1 NOT_1986 (.Y(g8858),.A(g8743));
INVX1 NOT_1987 (.Y(g4671),.A(g3354));
INVX1 NOT_1988 (.Y(g2880),.A(I6028));
INVX1 NOT_1989 (.Y(g4428),.A(I7776));
INVX1 NOT_1990 (.Y(g2537),.A(I5646));
INVX1 NOT_1991 (.Y(I10546),.A(g5914));
INVX1 NOT_1992 (.Y(g5896),.A(I9525));
INVX1 NOT_1993 (.Y(g4430),.A(I7782));
INVX1 NOT_1994 (.Y(I14546),.A(g9312));
INVX1 NOT_1995 (.Y(I7438),.A(g3461));
INVX1 NOT_1996 (.Y(g3164),.A(I6370));
INVX1 NOT_1997 (.Y(g3364),.A(g3121));
INVX1 NOT_1998 (.Y(I7009),.A(g2913));
INVX1 NOT_1999 (.Y(I10024),.A(g5700));
INVX1 NOT_2000 (.Y(I8204),.A(g3976));
INVX1 NOT_2001 (.Y(I12631),.A(g7705));
INVX1 NOT_2002 (.Y(g8115),.A(g7953));
INVX1 NOT_2003 (.Y(g4564),.A(g3880));
INVX1 NOT_2004 (.Y(g8251),.A(I13166));
INVX1 NOT_2005 (.Y(g8315),.A(I13329));
INVX1 NOT_2006 (.Y(g2612),.A(I5737));
INVX1 NOT_2007 (.Y(I15326),.A(g10025));
INVX1 NOT_2008 (.Y(g2017),.A(g1218));
INVX1 NOT_2009 (.Y(g6284),.A(I10111));
INVX1 NOT_2010 (.Y(g2243),.A(I5248));
INVX1 NOT_2011 (.Y(g8447),.A(I13639));
INVX1 NOT_2012 (.Y(I6580),.A(g3186));
INVX1 NOT_2013 (.Y(g3770),.A(I6985));
INVX1 NOT_2014 (.Y(g6239),.A(I9988));
INVX1 NOT_2015 (.Y(g10794),.A(I16496));
INVX1 NOT_2016 (.Y(I15536),.A(g10111));
INVX1 NOT_2017 (.Y(g10395),.A(g10320));
INVX1 NOT_2018 (.Y(g5419),.A(I8858));
INVX1 NOT_2019 (.Y(g9804),.A(I14939));
INVX1 NOT_2020 (.Y(g10262),.A(g10142));
INVX1 NOT_2021 (.Y(g7683),.A(g7148));
INVX1 NOT_2022 (.Y(g11040),.A(I16781));
INVX1 NOT_2023 (.Y(g10899),.A(g10803));
INVX1 NOT_2024 (.Y(g6591),.A(I10553));
INVX1 NOT_2025 (.Y(I11412),.A(g6411));
INVX1 NOT_2026 (.Y(g5052),.A(g4394));
INVX1 NOT_2027 (.Y(I13412),.A(g8142));
INVX1 NOT_2028 (.Y(I5101),.A(g1960));
INVX1 NOT_2029 (.Y(g8874),.A(I14194));
INVX1 NOT_2030 (.Y(g3532),.A(g3164));
INVX1 NOT_2031 (.Y(g7778),.A(I12499));
INVX1 NOT_2032 (.Y(g2234),.A(g87));
INVX1 NOT_2033 (.Y(g6853),.A(I10917));
INVX1 NOT_2034 (.Y(I10126),.A(g5682));
INVX1 NOT_2035 (.Y(I10659),.A(g6038));
INVX1 NOT_2036 (.Y(I16574),.A(g10821));
INVX1 NOT_2037 (.Y(g2629),.A(g2001));
INVX1 NOT_2038 (.Y(g4638),.A(g3354));
INVX1 NOT_2039 (.Y(g2328),.A(g1882));
INVX1 NOT_2040 (.Y(I12289),.A(g7142));
INVX1 NOT_2041 (.Y(I6968),.A(g2881));
INVX1 NOT_2042 (.Y(g6420),.A(I10334));
INVX1 NOT_2043 (.Y(g11621),.A(I17681));
INVX1 NOT_2044 (.Y(g2130),.A(I5057));
INVX1 NOT_2045 (.Y(g10191),.A(I15551));
INVX1 NOT_2046 (.Y(g2542),.A(g1868));
INVX1 NOT_2047 (.Y(I8973),.A(g4488));
INVX1 NOT_2048 (.Y(g2330),.A(g1891));
INVX1 NOT_2049 (.Y(g7735),.A(I12384));
INVX1 NOT_2050 (.Y(I16311),.A(g10584));
INVX1 NOT_2051 (.Y(g4308),.A(g3863));
INVX1 NOT_2052 (.Y(I11228),.A(g6471));
INVX1 NOT_2053 (.Y(I17231),.A(g11303));
INVX1 NOT_2054 (.Y(g7782),.A(I12511));
INVX1 NOT_2055 (.Y(g6559),.A(g5758));
INVX1 NOT_2056 (.Y(I12571),.A(g7509));
INVX1 NOT_2057 (.Y(g3012),.A(I6247));
INVX1 NOT_2058 (.Y(I11011),.A(g6340));
INVX1 NOT_2059 (.Y(I5751),.A(g2296));
INVX1 NOT_2060 (.Y(g8595),.A(I13840));
INVX1 NOT_2061 (.Y(g6931),.A(I11055));
INVX1 NOT_2062 (.Y(g5728),.A(I9276));
INVX1 NOT_2063 (.Y(g5486),.A(g4395));
INVX1 NOT_2064 (.Y(I10296),.A(g6242));
INVX1 NOT_2065 (.Y(I11716),.A(g7026));
INVX1 NOT_2066 (.Y(g5730),.A(I9282));
INVX1 NOT_2067 (.Y(g5504),.A(g4419));
INVX1 NOT_2068 (.Y(g7949),.A(g7422));
INVX1 NOT_2069 (.Y(g4217),.A(I7468));
INVX1 NOT_2070 (.Y(g11183),.A(I16950));
INVX1 NOT_2071 (.Y(I8123),.A(g3630));
INVX1 NOT_2072 (.Y(g3990),.A(g3121));
INVX1 NOT_2073 (.Y(g2554),.A(I5672));
INVX1 NOT_2074 (.Y(g4758),.A(g3586));
INVX1 NOT_2075 (.Y(g4066),.A(I7191));
INVX1 NOT_2076 (.Y(g8272),.A(I13188));
INVX1 NOT_2077 (.Y(I16592),.A(g10781));
INVX1 NOT_2078 (.Y(g4589),.A(I7996));
INVX1 NOT_2079 (.Y(g5185),.A(g4682));
INVX1 NOT_2080 (.Y(g11397),.A(I17234));
INVX1 NOT_2081 (.Y(g5881),.A(g5361));
INVX1 NOT_2082 (.Y(g7627),.A(I12223));
INVX1 NOT_2083 (.Y(g9094),.A(g8892));
INVX1 NOT_2084 (.Y(I5041),.A(g1179));
INVX1 NOT_2085 (.Y(I9135),.A(g5198));
INVX1 NOT_2086 (.Y(g4466),.A(I7833));
INVX1 NOT_2087 (.Y(g1992),.A(g782));
INVX1 NOT_2088 (.Y(g6905),.A(I11011));
INVX1 NOT_2089 (.Y(g8978),.A(I14355));
INVX1 NOT_2090 (.Y(I5441),.A(g919));
INVX1 NOT_2091 (.Y(g3371),.A(g2837));
INVX1 NOT_2092 (.Y(g11062),.A(g10937));
INVX1 NOT_2093 (.Y(I10060),.A(g5752));
INVX1 NOT_2094 (.Y(g2213),.A(g1110));
INVX1 NOT_2095 (.Y(g11509),.A(I17546));
INVX1 NOT_2096 (.Y(g7998),.A(I12822));
INVX1 NOT_2097 (.Y(g10247),.A(I15639));
INVX1 NOT_2098 (.Y(g4165),.A(g3164));
INVX1 NOT_2099 (.Y(g4365),.A(g3880));
INVX1 NOT_2100 (.Y(I13627),.A(g8326));
INVX1 NOT_2101 (.Y(g5425),.A(g4300));
INVX1 NOT_2102 (.Y(g10389),.A(g10307));
INVX1 NOT_2103 (.Y(g10926),.A(g10827));
INVX1 NOT_2104 (.Y(I10855),.A(g6685));
INVX1 NOT_2105 (.Y(I13959),.A(g8451));
INVX1 NOT_2106 (.Y(I13379),.A(g8133));
INVX1 NOT_2107 (.Y(g11508),.A(I17543));
INVX1 NOT_2108 (.Y(g4711),.A(I8061));
INVX1 NOT_2109 (.Y(g6100),.A(I9759));
INVX1 NOT_2110 (.Y(I11112),.A(g6445));
INVX1 NOT_2111 (.Y(g8982),.A(I14367));
INVX1 NOT_2112 (.Y(g11634),.A(I17716));
INVX1 NOT_2113 (.Y(g10612),.A(I16286));
INVX1 NOT_2114 (.Y(g6300),.A(I10159));
INVX1 NOT_2115 (.Y(g7603),.A(I12159));
INVX1 NOT_2116 (.Y(g4055),.A(g3144));
INVX1 NOT_2117 (.Y(g7039),.A(I11204));
INVX1 NOT_2118 (.Y(I9749),.A(g5266));
INVX1 NOT_2119 (.Y(g10388),.A(g10305));
INVX1 NOT_2120 (.Y(I8351),.A(g4794));
INVX1 NOT_2121 (.Y(g8234),.A(g7826));
INVX1 NOT_2122 (.Y(g2902),.A(I6061));
INVX1 NOT_2123 (.Y(g7439),.A(I11833));
INVX1 NOT_2124 (.Y(g8128),.A(I12993));
INVX1 NOT_2125 (.Y(g8328),.A(I13364));
INVX1 NOT_2126 (.Y(g7850),.A(I12647));
INVX1 NOT_2127 (.Y(g10534),.A(I16169));
INVX1 NOT_2128 (.Y(g10098),.A(I15332));
INVX1 NOT_2129 (.Y(I17456),.A(g11453));
INVX1 NOT_2130 (.Y(g4333),.A(g4144));
INVX1 NOT_2131 (.Y(I7837),.A(g4158));
INVX1 NOT_2132 (.Y(g8330),.A(I13370));
INVX1 NOT_2133 (.Y(g10251),.A(g10195));
INVX1 NOT_2134 (.Y(g10272),.A(g10168));
INVX1 NOT_2135 (.Y(g2090),.A(I4920));
INVX1 NOT_2136 (.Y(g4774),.A(I8136));
INVX1 NOT_2137 (.Y(I7462),.A(g3721));
INVX1 NOT_2138 (.Y(I9798),.A(g5415));
INVX1 NOT_2139 (.Y(I13096),.A(g7925));
INVX1 NOT_2140 (.Y(g2166),.A(I5101));
INVX1 NOT_2141 (.Y(g6750),.A(I10759));
INVX1 NOT_2142 (.Y(g9264),.A(I14477));
INVX1 NOT_2143 (.Y(I6424),.A(g2462));
INVX1 NOT_2144 (.Y(g7702),.A(g7079));
INVX1 NOT_2145 (.Y(g4196),.A(I7405));
INVX1 NOT_2146 (.Y(g5678),.A(I9191));
INVX1 NOT_2147 (.Y(I10503),.A(g5858));
INVX1 NOT_2148 (.Y(I16413),.A(g10663));
INVX1 NOT_2149 (.Y(g10462),.A(I15977));
INVX1 NOT_2150 (.Y(g4396),.A(I7735));
INVX1 NOT_2151 (.Y(g3138),.A(I6356));
INVX1 NOT_2152 (.Y(g8800),.A(I14123));
INVX1 NOT_2153 (.Y(I14503),.A(g8920));
INVX1 NOT_2154 (.Y(I8410),.A(g4283));
INVX1 NOT_2155 (.Y(g2056),.A(I4859));
INVX1 NOT_2156 (.Y(I16691),.A(g10788));
INVX1 NOT_2157 (.Y(g9360),.A(I14579));
INVX1 NOT_2158 (.Y(g3109),.A(g2482));
INVX1 NOT_2159 (.Y(g3791),.A(I7014));
INVX1 NOT_2160 (.Y(g2456),.A(g1397));
INVX1 NOT_2161 (.Y(g7919),.A(g7512));
INVX1 NOT_2162 (.Y(g10032),.A(I15232));
INVX1 NOT_2163 (.Y(g2529),.A(I5638));
INVX1 NOT_2164 (.Y(g2649),.A(g2005));
INVX1 NOT_2165 (.Y(g10140),.A(I15418));
INVX1 NOT_2166 (.Y(g4780),.A(g3440));
INVX1 NOT_2167 (.Y(I8839),.A(g4484));
INVX1 NOT_2168 (.Y(g6040),.A(I9655));
INVX1 NOT_2169 (.Y(g2348),.A(I5418));
INVX1 NOT_2170 (.Y(I6077),.A(g2349));
INVX1 NOT_2171 (.Y(g11574),.A(g11561));
INVX1 NOT_2172 (.Y(g11452),.A(I17413));
INVX1 NOT_2173 (.Y(g11047),.A(I16802));
INVX1 NOT_2174 (.Y(g5682),.A(I9199));
INVX1 NOT_2175 (.Y(g5766),.A(I9346));
INVX1 NOT_2176 (.Y(g5105),.A(I8487));
INVX1 NOT_2177 (.Y(g4509),.A(I7906));
INVX1 NOT_2178 (.Y(g6440),.A(g6150));
INVX1 NOT_2179 (.Y(g1976),.A(g643));
INVX1 NOT_2180 (.Y(g11205),.A(g11112));
INVX1 NOT_2181 (.Y(I6477),.A(g2069));
INVX1 NOT_2182 (.Y(I9632),.A(g5557));
INVX1 NOT_2183 (.Y(g7952),.A(g7427));
INVX1 NOT_2184 (.Y(I15311),.A(g10013));
INVX1 NOT_2185 (.Y(g9450),.A(g9097));
INVX1 NOT_2186 (.Y(g5305),.A(g4378));
INVX1 NOT_2187 (.Y(g5801),.A(g5320));
INVX1 NOT_2188 (.Y(I5734),.A(g2097));
INVX1 NOT_2189 (.Y(I6523),.A(g2819));
INVX1 NOT_2190 (.Y(g2155),.A(I5070));
INVX1 NOT_2191 (.Y(I4820),.A(g865));
INVX1 NOT_2192 (.Y(I17243),.A(g11396));
INVX1 NOT_2193 (.Y(g2355),.A(I5435));
INVX1 NOT_2194 (.Y(g2851),.A(I5979));
INVX1 NOT_2195 (.Y(I7249),.A(g2833));
INVX1 NOT_2196 (.Y(I12559),.A(g7477));
INVX1 NOT_2197 (.Y(I14315),.A(g8815));
INVX1 NOT_2198 (.Y(I6643),.A(g3008));
INVX1 NOT_2199 (.Y(g8213),.A(g7826));
INVX1 NOT_2200 (.Y(I10819),.A(g6706));
INVX1 NOT_2201 (.Y(g11311),.A(I17100));
INVX1 NOT_2202 (.Y(I10910),.A(g6703));
INVX1 NOT_2203 (.Y(I12424),.A(g7635));
INVX1 NOT_2204 (.Y(I9102),.A(g5586));
INVX1 NOT_2205 (.Y(I9208),.A(g5047));
INVX1 NOT_2206 (.Y(g3707),.A(g2920));
INVX1 NOT_2207 (.Y(I9302),.A(g5576));
INVX1 NOT_2208 (.Y(I14910),.A(g9532));
INVX1 NOT_2209 (.Y(g7616),.A(I12196));
INVX1 NOT_2210 (.Y(g7561),.A(I12015));
INVX1 NOT_2211 (.Y(g4067),.A(I7194));
INVX1 NOT_2212 (.Y(g3759),.A(I6958));
INVX1 NOT_2213 (.Y(I8278),.A(g4495));
INVX1 NOT_2214 (.Y(I14257),.A(g8805));
INVX1 NOT_2215 (.Y(g5748),.A(I9320));
INVX1 NOT_2216 (.Y(I10979),.A(g6565));
INVX1 NOT_2217 (.Y(g2964),.A(I6193));
INVX1 NOT_2218 (.Y(g4418),.A(I7760));
INVX1 NOT_2219 (.Y(I9869),.A(g5405));
INVX1 NOT_2220 (.Y(g4467),.A(g3829));
INVX1 NOT_2221 (.Y(I15072),.A(g9713));
INVX1 NOT_2222 (.Y(I14979),.A(g9671));
INVX1 NOT_2223 (.Y(g4290),.A(g3586));
INVX1 NOT_2224 (.Y(I10111),.A(g5754));
INVX1 NOT_2225 (.Y(I14055),.A(g8650));
INVX1 NOT_2226 (.Y(g10871),.A(I16583));
INVX1 NOT_2227 (.Y(g11051),.A(I16814));
INVX1 NOT_2228 (.Y(I5992),.A(g2195));
INVX1 NOT_2229 (.Y(g7004),.A(I11143));
INVX1 NOT_2230 (.Y(I16583),.A(g10848));
INVX1 NOT_2231 (.Y(g11072),.A(g10913));
INVX1 NOT_2232 (.Y(I17773),.A(g11650));
INVX1 NOT_2233 (.Y(I15592),.A(g10163));
INVX1 NOT_2234 (.Y(I15756),.A(g10266));
INVX1 NOT_2235 (.Y(g7527),.A(g7148));
INVX1 NOT_2236 (.Y(I17268),.A(g11351));
INVX1 NOT_2237 (.Y(I6742),.A(g3326));
INVX1 NOT_2238 (.Y(I12544),.A(g7669));
INVX1 NOT_2239 (.Y(g4093),.A(g2965));
INVX1 NOT_2240 (.Y(I8282),.A(g4770));
INVX1 NOT_2241 (.Y(g6151),.A(I9872));
INVX1 NOT_2242 (.Y(g7764),.A(I12457));
INVX1 NOT_2243 (.Y(g4256),.A(g3664));
INVX1 NOT_2244 (.Y(g6648),.A(I10607));
INVX1 NOT_2245 (.Y(g9777),.A(g9474));
INVX1 NOT_2246 (.Y(g7546),.A(I11970));
INVX1 NOT_2247 (.Y(I5080),.A(g36));
INVX1 NOT_2248 (.Y(I15350),.A(g10001));
INVX1 NOT_2249 (.Y(I10384),.A(g5842));
INVX1 NOT_2250 (.Y(g10162),.A(I15482));
INVX1 NOT_2251 (.Y(g3715),.A(g2920));
INVX1 NOT_2252 (.Y(I9265),.A(g5085));
INVX1 NOT_2253 (.Y(I16787),.A(g10896));
INVX1 NOT_2254 (.Y(g11350),.A(g11287));
INVX1 NOT_2255 (.Y(I5713),.A(g2436));
INVX1 NOT_2256 (.Y(I15820),.A(g10204));
INVX1 NOT_2257 (.Y(g5091),.A(g4385));
INVX1 NOT_2258 (.Y(g8056),.A(g7671));
INVX1 NOT_2259 (.Y(I13317),.A(g8093));
INVX1 NOT_2260 (.Y(I12610),.A(g7627));
INVX1 NOT_2261 (.Y(g4181),.A(I7360));
INVX1 NOT_2262 (.Y(I6754),.A(g2906));
INVX1 NOT_2263 (.Y(g8529),.A(I13738));
INVX1 NOT_2264 (.Y(I14094),.A(g8700));
INVX1 NOT_2265 (.Y(g4381),.A(g3914));
INVX1 NOT_2266 (.Y(g7925),.A(g7476));
INVX1 NOT_2267 (.Y(I9786),.A(g5396));
INVX1 NOT_2268 (.Y(g2118),.A(g1854));
INVX1 NOT_2269 (.Y(g8348),.A(I13424));
INVX1 NOT_2270 (.Y(I12255),.A(g7203));
INVX1 NOT_2271 (.Y(I6273),.A(g2482));
INVX1 NOT_2272 (.Y(g2872),.A(I6016));
INVX1 NOT_2273 (.Y(I16105),.A(g10382));
INVX1 NOT_2274 (.Y(g10629),.A(g10583));
INVX1 NOT_2275 (.Y(I10150),.A(g5705));
INVX1 NOT_2276 (.Y(g5169),.A(g4596));
INVX1 NOT_2277 (.Y(g4197),.A(I7408));
INVX1 NOT_2278 (.Y(I10801),.A(g6536));
INVX1 NOT_2279 (.Y(g8155),.A(I13048));
INVX1 NOT_2280 (.Y(g11396),.A(I17231));
INVX1 NOT_2281 (.Y(I13002),.A(g8045));
INVX1 NOT_2282 (.Y(g8355),.A(I13445));
INVX1 NOT_2283 (.Y(g10220),.A(I15592));
INVX1 NOT_2284 (.Y(g5007),.A(I8379));
INVX1 NOT_2285 (.Y(I13057),.A(g7843));
INVX1 NOT_2286 (.Y(g2652),.A(g2008));
INVX1 NOT_2287 (.Y(g2057),.A(g754));
INVX1 NOT_2288 (.Y(g10628),.A(I16307));
INVX1 NOT_2289 (.Y(I12678),.A(g7376));
INVX1 NOT_2290 (.Y(I13128),.A(g7976));
INVX1 NOT_2291 (.Y(g2843),.A(I5963));
INVX1 NOT_2292 (.Y(g10911),.A(I16685));
INVX1 NOT_2293 (.Y(g7320),.A(I11608));
INVX1 NOT_2294 (.Y(g2989),.A(g2135));
INVX1 NOT_2295 (.Y(g3539),.A(g3015));
INVX1 NOT_2296 (.Y(g4263),.A(g3586));
INVX1 NOT_2297 (.Y(I13245),.A(g8269));
INVX1 NOT_2298 (.Y(I11626),.A(g7042));
INVX1 NOT_2299 (.Y(I16769),.A(g10894));
INVX1 NOT_2300 (.Y(g5718),.A(I9256));
INVX1 NOT_2301 (.Y(I12460),.A(g7569));
INVX1 NOT_2302 (.Y(I12939),.A(g7977));
INVX1 NOT_2303 (.Y(g5767),.A(I9349));
INVX1 NOT_2304 (.Y(I15691),.A(g10233));
INVX1 NOT_2305 (.Y(I9296),.A(g4908));
INVX1 NOT_2306 (.Y(I10018),.A(g5862));
INVX1 NOT_2307 (.Y(I11299),.A(g6727));
INVX1 NOT_2308 (.Y(I13323),.A(g8203));
INVX1 NOT_2309 (.Y(I7176),.A(g2623));
INVX1 NOT_2310 (.Y(I5976),.A(g2186));
INVX1 NOT_2311 (.Y(g2549),.A(g1386));
INVX1 NOT_2312 (.Y(I6572),.A(g2853));
INVX1 NOT_2313 (.Y(I10526),.A(g6161));
INVX1 NOT_2314 (.Y(g8063),.A(I12907));
INVX1 NOT_2315 (.Y(g2834),.A(I5952));
INVX1 NOT_2316 (.Y(g2971),.A(g2046));
INVX1 NOT_2317 (.Y(g6172),.A(I9901));
INVX1 NOT_2318 (.Y(g6278),.A(I10093));
INVX1 NOT_2319 (.Y(g7617),.A(I12199));
INVX1 NOT_2320 (.Y(I7405),.A(g3861));
INVX1 NOT_2321 (.Y(g7906),.A(I12694));
INVX1 NOT_2322 (.Y(g7789),.A(I12532));
INVX1 NOT_2323 (.Y(g11405),.A(I17258));
INVX1 NOT_2324 (.Y(g5261),.A(g4640));
INVX1 NOT_2325 (.Y(g10591),.A(I16258));
INVX1 NOT_2326 (.Y(I6543),.A(g3186));
INVX1 NOT_2327 (.Y(g3362),.A(I6546));
INVX1 NOT_2328 (.Y(g3419),.A(g3104));
INVX1 NOT_2329 (.Y(I7829),.A(g3425));
INVX1 NOT_2330 (.Y(g6667),.A(I10630));
INVX1 NOT_2331 (.Y(g7516),.A(g7148));
INVX1 NOT_2332 (.Y(g4562),.A(I7973));
INVX1 NOT_2333 (.Y(g6343),.A(I10248));
INVX1 NOT_2334 (.Y(g10754),.A(I16439));
INVX1 NOT_2335 (.Y(g9353),.A(I14564));
INVX1 NOT_2336 (.Y(g3052),.A(I6264));
INVX1 NOT_2337 (.Y(g10355),.A(I15829));
INVX1 NOT_2338 (.Y(g5415),.A(I8848));
INVX1 NOT_2339 (.Y(g6282),.A(I10105));
INVX1 NOT_2340 (.Y(g7771),.A(I12478));
INVX1 NOT_2341 (.Y(g6566),.A(g5791));
INVX1 NOT_2342 (.Y(I11737),.A(g7027));
INVX1 NOT_2343 (.Y(g8279),.A(I13209));
INVX1 NOT_2344 (.Y(g2121),.A(I5041));
INVX1 NOT_2345 (.Y(g4631),.A(g3820));
INVX1 NOT_2346 (.Y(I12875),.A(g7638));
INVX1 NOT_2347 (.Y(g10825),.A(I16537));
INVX1 NOT_2348 (.Y(I10917),.A(g6732));
INVX1 NOT_2349 (.Y(I15583),.A(g10157));
INVX1 NOT_2350 (.Y(g9802),.A(g9490));
INVX1 NOT_2351 (.Y(g1999),.A(g806));
INVX1 NOT_2352 (.Y(I11232),.A(g6537));
INVX1 NOT_2353 (.Y(g4257),.A(g3664));
INVX1 NOT_2354 (.Y(g6134),.A(I9839));
INVX1 NOT_2355 (.Y(g5664),.A(I9153));
INVX1 NOT_2356 (.Y(g8318),.A(I13338));
INVX1 NOT_2357 (.Y(g8872),.A(I14188));
INVX1 NOT_2358 (.Y(I9706),.A(g5221));
INVX1 NOT_2359 (.Y(g2232),.A(I5221));
INVX1 NOT_2360 (.Y(g10172),.A(I15510));
INVX1 NOT_2361 (.Y(g11046),.A(I16799));
INVX1 NOT_2362 (.Y(g3086),.A(g2276));
INVX1 NOT_2363 (.Y(g5203),.A(g4640));
INVX1 NOT_2364 (.Y(g2253),.A(g100));
INVX1 NOT_2365 (.Y(g3728),.A(I6904));
INVX1 NOT_2366 (.Y(g2813),.A(I5913));
INVX1 NOT_2367 (.Y(I9029),.A(g4781));
INVX1 NOT_2368 (.Y(g8989),.A(I14388));
INVX1 NOT_2369 (.Y(I14077),.A(g8758));
INVX1 NOT_2370 (.Y(I9171),.A(g4902));
INVX1 NOT_2371 (.Y(g6555),.A(g5740));
INVX1 NOT_2372 (.Y(I10706),.A(g6080));
INVX1 NOT_2373 (.Y(I9371),.A(g5075));
INVX1 NOT_2374 (.Y(g6804),.A(I10822));
INVX1 NOT_2375 (.Y(I15787),.A(g10269));
INVX1 NOT_2376 (.Y(I6414),.A(g2342));
INVX1 NOT_2377 (.Y(g3730),.A(g3015));
INVX1 NOT_2378 (.Y(g2909),.A(I6080));
INVX1 NOT_2379 (.Y(I9956),.A(g5485));
INVX1 NOT_2380 (.Y(I10689),.A(g6059));
INVX1 NOT_2381 (.Y(g3385),.A(g3121));
INVX1 NOT_2382 (.Y(I5383),.A(g886));
INVX1 NOT_2383 (.Y(I15302),.A(g10007));
INVX1 NOT_2384 (.Y(g11357),.A(I17182));
INVX1 NOT_2385 (.Y(g7991),.A(I12809));
INVX1 NOT_2386 (.Y(I6513),.A(g2812));
INVX1 NOT_2387 (.Y(g2606),.A(I5719));
INVX1 NOT_2388 (.Y(g10319),.A(g10270));
INVX1 NOT_2389 (.Y(g4441),.A(g3914));
INVX1 NOT_2390 (.Y(g6113),.A(I9792));
INVX1 NOT_2391 (.Y(g6313),.A(I10198));
INVX1 NOT_2392 (.Y(g7078),.A(I11309));
INVX1 NOT_2393 (.Y(g7340),.A(I11668));
INVX1 NOT_2394 (.Y(I10102),.A(g5730));
INVX1 NOT_2395 (.Y(I16778),.A(g10891));
INVX1 NOT_2396 (.Y(I13831),.A(g8560));
INVX1 NOT_2397 (.Y(g10318),.A(I15752));
INVX1 NOT_2398 (.Y(I8050),.A(g4089));
INVX1 NOT_2399 (.Y(I13445),.A(g8149));
INVX1 NOT_2400 (.Y(I5588),.A(g1203));
INVX1 NOT_2401 (.Y(g8121),.A(I12978));
INVX1 NOT_2402 (.Y(g10227),.A(I15601));
INVX1 NOT_2403 (.Y(g7907),.A(g7664));
INVX1 NOT_2404 (.Y(I6436),.A(g2351));
INVX1 NOT_2405 (.Y(I6679),.A(g2902));
INVX1 NOT_2406 (.Y(g8321),.A(I13347));
INVX1 NOT_2407 (.Y(g4673),.A(g4013));
INVX1 NOT_2408 (.Y(g6202),.A(g5426));
INVX1 NOT_2409 (.Y(g8670),.A(g8551));
INVX1 NOT_2410 (.Y(g5689),.A(I9216));
INVX1 NOT_2411 (.Y(I8996),.A(g4757));
INVX1 NOT_2412 (.Y(I9684),.A(g5426));
INVX1 NOT_2413 (.Y(g7035),.A(I11194));
INVX1 NOT_2414 (.Y(I15768),.A(g10249));
INVX1 NOT_2415 (.Y(I9138),.A(g5210));
INVX1 NOT_2416 (.Y(I9639),.A(g5126));
INVX1 NOT_2417 (.Y(g7959),.A(I12751));
INVX1 NOT_2418 (.Y(I10066),.A(g5778));
INVX1 NOT_2419 (.Y(I9338),.A(g5576));
INVX1 NOT_2420 (.Y(I10231),.A(g6111));
INVX1 NOT_2421 (.Y(g8625),.A(g8487));
INVX1 NOT_2422 (.Y(g7082),.A(I11315));
INVX1 NOT_2423 (.Y(g2586),.A(g1972));
INVX1 NOT_2424 (.Y(g5216),.A(g4445));
INVX1 NOT_2425 (.Y(g10540),.A(I16187));
INVX1 NOT_2426 (.Y(I17410),.A(g11419));
INVX1 NOT_2427 (.Y(g6094),.A(I9749));
INVX1 NOT_2428 (.Y(I11498),.A(g6578));
INVX1 NOT_2429 (.Y(I12595),.A(g7706));
INVX1 NOT_2430 (.Y(I16647),.A(g10866));
INVX1 NOT_2431 (.Y(g10058),.A(I15281));
INVX1 NOT_2432 (.Y(I16356),.A(g10597));
INVX1 NOT_2433 (.Y(g4669),.A(g4013));
INVX1 NOT_2434 (.Y(I8724),.A(g4791));
INVX1 NOT_2435 (.Y(g6567),.A(I10495));
INVX1 NOT_2436 (.Y(g5671),.A(I9174));
INVX1 NOT_2437 (.Y(g4368),.A(I7665));
INVX1 NOT_2438 (.Y(I11989),.A(g6919));
INVX1 NOT_2439 (.Y(I17666),.A(g11603));
INVX1 NOT_2440 (.Y(I10885),.A(g6332));
INVX1 NOT_2441 (.Y(I8379),.A(g4231));
INVX1 NOT_2442 (.Y(g3331),.A(I6510));
INVX1 NOT_2443 (.Y(g10203),.A(g10177));
INVX1 NOT_2444 (.Y(I14876),.A(g9526));
INVX1 NOT_2445 (.Y(I11611),.A(g6913));
INVX1 NOT_2446 (.Y(g7656),.A(I12265));
INVX1 NOT_2447 (.Y(g4772),.A(g3440));
INVX1 NOT_2448 (.Y(g3406),.A(I6611));
INVX1 NOT_2449 (.Y(I11722),.A(g7034));
INVX1 NOT_2450 (.Y(I7399),.A(g4113));
INVX1 NOT_2451 (.Y(g10044),.A(I15263));
INVX1 NOT_2452 (.Y(g3635),.A(I6812));
INVX1 NOT_2453 (.Y(I6022),.A(g2258));
INVX1 NOT_2454 (.Y(g4458),.A(I7817));
INVX1 NOT_2455 (.Y(g2570),.A(g207));
INVX1 NOT_2456 (.Y(g2860),.A(I5998));
INVX1 NOT_2457 (.Y(g2341),.A(I5403));
INVX1 NOT_2458 (.Y(g9262),.A(I14473));
INVX1 NOT_2459 (.Y(g3682),.A(g2920));
INVX1 NOT_2460 (.Y(g6593),.A(I10557));
INVX1 NOT_2461 (.Y(I9759),.A(g5344));
INVX1 NOT_2462 (.Y(g8519),.A(I13726));
INVX1 NOT_2463 (.Y(g3105),.A(g2482));
INVX1 NOT_2464 (.Y(g7915),.A(g7473));
INVX1 NOT_2465 (.Y(g3305),.A(I6474));
INVX1 NOT_2466 (.Y(g10281),.A(g10162));
INVX1 NOT_2467 (.Y(g98),.A(I4783));
INVX1 NOT_2468 (.Y(g2645),.A(g1991));
INVX1 NOT_2469 (.Y(I8835),.A(g4791));
INVX1 NOT_2470 (.Y(g5826),.A(I9440));
INVX1 NOT_2471 (.Y(I12418),.A(g7568));
INVX1 NOT_2472 (.Y(I12822),.A(g7677));
INVX1 NOT_2473 (.Y(g10902),.A(I16660));
INVX1 NOT_2474 (.Y(g10377),.A(I15855));
INVX1 NOT_2475 (.Y(g8606),.A(g8481));
INVX1 NOT_2476 (.Y(g7214),.A(I11450));
INVX1 NOT_2477 (.Y(I6947),.A(g2860));
INVX1 NOT_2478 (.Y(g10120),.A(I15368));
INVX1 NOT_2479 (.Y(g4011),.A(I7151));
INVX1 NOT_2480 (.Y(g9076),.A(g8892));
INVX1 NOT_2481 (.Y(g5741),.A(I9305));
INVX1 NOT_2482 (.Y(g3748),.A(g2971));
INVX1 NOT_2483 (.Y(g4411),.A(I7743));
INVX1 NOT_2484 (.Y(g4734),.A(g3586));
INVX1 NOT_2485 (.Y(I11342),.A(g6686));
INVX1 NOT_2486 (.Y(g9889),.A(I15072));
INVX1 NOT_2487 (.Y(g7110),.A(I11345));
INVX1 NOT_2488 (.Y(g6264),.A(I10051));
INVX1 NOT_2489 (.Y(g7310),.A(I11578));
INVX1 NOT_2490 (.Y(I6560),.A(g2845));
INVX1 NOT_2491 (.Y(I7291),.A(g3212));
INVX1 NOT_2492 (.Y(I8611),.A(g4562));
INVX1 NOT_2493 (.Y(I10456),.A(g5844));
INVX1 NOT_2494 (.Y(I15482),.A(g10115));
INVX1 NOT_2495 (.Y(g5638),.A(I9077));
INVX1 NOT_2496 (.Y(g3226),.A(I6403));
INVX1 NOT_2497 (.Y(g6933),.A(I11061));
INVX1 NOT_2498 (.Y(g7663),.A(I12282));
INVX1 NOT_2499 (.Y(I11650),.A(g6938));
INVX1 NOT_2500 (.Y(g10699),.A(I16376));
INVX1 NOT_2501 (.Y(g2607),.A(I5722));
INVX1 NOT_2502 (.Y(I12853),.A(g7638));
INVX1 NOT_2503 (.Y(I16897),.A(g10947));
INVX1 NOT_2504 (.Y(I5240),.A(g64));
INVX1 NOT_2505 (.Y(g2962),.A(I6183));
INVX1 NOT_2506 (.Y(g6521),.A(I10437));
INVX1 NOT_2507 (.Y(I17084),.A(g11249));
INVX1 NOT_2508 (.Y(g4474),.A(g3820));
INVX1 NOT_2509 (.Y(g10290),.A(I15694));
INVX1 NOT_2510 (.Y(g2158),.A(I5077));
INVX1 NOT_2511 (.Y(g6050),.A(I9677));
INVX1 NOT_2512 (.Y(g6641),.A(I10598));
INVX1 NOT_2513 (.Y(I11198),.A(g6521));
INVX1 NOT_2514 (.Y(I9498),.A(g5081));
INVX1 NOT_2515 (.Y(I12589),.A(g7571));
INVX1 NOT_2516 (.Y(g10698),.A(I16373));
INVX1 NOT_2517 (.Y(g2506),.A(g636));
INVX1 NOT_2518 (.Y(g6450),.A(I10378));
INVX1 NOT_2519 (.Y(I6037),.A(g2560));
INVX1 NOT_2520 (.Y(I17321),.A(g11348));
INVX1 NOT_2521 (.Y(g5883),.A(g5309));
INVX1 NOT_2522 (.Y(I10314),.A(g6251));
INVX1 NOT_2523 (.Y(g7402),.A(g6860));
INVX1 NOT_2524 (.Y(I6495),.A(g2076));
INVX1 NOT_2525 (.Y(I9833),.A(g5197));
INVX1 NOT_2526 (.Y(I17179),.A(g11307));
INVX1 NOT_2527 (.Y(I11528),.A(g6796));
INVX1 NOT_2528 (.Y(I6102),.A(g2240));
INVX1 NOT_2529 (.Y(I16717),.A(g10779));
INVX1 NOT_2530 (.Y(I17531),.A(g11488));
INVX1 NOT_2531 (.Y(I7694),.A(g3742));
INVX1 NOT_2532 (.Y(I11330),.A(g6571));
INVX1 NOT_2533 (.Y(I6302),.A(g2243));
INVX1 NOT_2534 (.Y(g3373),.A(I6565));
INVX1 NOT_2535 (.Y(I15778),.A(g10255));
INVX1 NOT_2536 (.Y(g7762),.A(I12451));
INVX1 NOT_2537 (.Y(g3491),.A(g2669));
INVX1 NOT_2538 (.Y(g4080),.A(g2903));
INVX1 NOT_2539 (.Y(I5116),.A(g40));
INVX1 NOT_2540 (.Y(g11081),.A(I16856));
INVX1 NOT_2541 (.Y(I7852),.A(g3438));
INVX1 NOT_2542 (.Y(I7923),.A(g3394));
INVX1 NOT_2543 (.Y(g5758),.A(I9338));
INVX1 NOT_2544 (.Y(g8141),.A(I13020));
INVX1 NOT_2545 (.Y(g8570),.A(I13803));
INVX1 NOT_2546 (.Y(g5066),.A(I8436));
INVX1 NOT_2547 (.Y(g5589),.A(I9001));
INVX1 NOT_2548 (.Y(g6724),.A(I10719));
INVX1 NOT_2549 (.Y(g8341),.A(I13403));
INVX1 NOT_2550 (.Y(I10054),.A(g5728));
INVX1 NOT_2551 (.Y(g2275),.A(g757));
INVX1 NOT_2552 (.Y(I9539),.A(g5354));
INVX1 NOT_2553 (.Y(I9896),.A(g5295));
INVX1 NOT_2554 (.Y(g4713),.A(g3546));
INVX1 NOT_2555 (.Y(I10243),.A(g5918));
INVX1 NOT_2556 (.Y(I11132),.A(g6451));
INVX1 NOT_2557 (.Y(I11869),.A(g6894));
INVX1 NOT_2558 (.Y(g7877),.A(g7479));
INVX1 NOT_2559 (.Y(I7701),.A(g3513));
INVX1 NOT_2560 (.Y(g3369),.A(I6557));
INVX1 NOT_2561 (.Y(I5565),.A(g1713));
INVX1 NOT_2562 (.Y(g3007),.A(I6240));
INVX1 NOT_2563 (.Y(g9339),.A(I14522));
INVX1 NOT_2564 (.Y(I15356),.A(g10013));
INVX1 NOT_2565 (.Y(g7657),.A(I12268));
INVX1 NOT_2566 (.Y(g6878),.A(I10966));
INVX1 NOT_2567 (.Y(I15826),.A(g10205));
INVX1 NOT_2568 (.Y(I6917),.A(g2832));
INVX1 NOT_2569 (.Y(I15380),.A(g10098));
INVX1 NOT_2570 (.Y(I4894),.A(g258));
INVX1 NOT_2571 (.Y(g2174),.A(g31));
INVX1 NOT_2572 (.Y(g3459),.A(I6661));
INVX1 NOT_2573 (.Y(g6289),.A(I10126));
INVX1 NOT_2574 (.Y(g9024),.A(I14409));
INVX1 NOT_2575 (.Y(g2374),.A(g591));
INVX1 NOT_2576 (.Y(I12616),.A(g7534));
INVX1 NOT_2577 (.Y(I9162),.A(g5035));
INVX1 NOT_2578 (.Y(g7556),.A(I11992));
INVX1 NOT_2579 (.Y(I9268),.A(g5305));
INVX1 NOT_2580 (.Y(I16723),.A(g10851));
INVX1 NOT_2581 (.Y(g3767),.A(I6976));
INVX1 NOT_2582 (.Y(g10547),.A(I16206));
INVX1 NOT_2583 (.Y(g9424),.A(g9076));
INVX1 NOT_2584 (.Y(g10895),.A(I16647));
INVX1 NOT_2585 (.Y(I7886),.A(g4076));
INVX1 NOT_2586 (.Y(I9362),.A(g5013));
INVX1 NOT_2587 (.Y(g6835),.A(I10885));
INVX1 NOT_2588 (.Y(g2985),.A(I6217));
INVX1 NOT_2589 (.Y(g9809),.A(I14944));
INVX1 NOT_2590 (.Y(g5827),.A(I9443));
INVX1 NOT_2591 (.Y(g6882),.A(I10974));
INVX1 NOT_2592 (.Y(g7928),.A(g7508));
INVX1 NOT_2593 (.Y(I10156),.A(g6100));
INVX1 NOT_2594 (.Y(I10655),.A(g6036));
INVX1 NOT_2595 (.Y(I15672),.A(g10132));
INVX1 NOT_2596 (.Y(g3582),.A(g3164));
INVX1 NOT_2597 (.Y(I16387),.A(g10629));
INVX1 NOT_2598 (.Y(I17334),.A(g11360));
INVX1 NOT_2599 (.Y(g6271),.A(I10072));
INVX1 NOT_2600 (.Y(I11225),.A(g6534));
INVX1 NOT_2601 (.Y(g10226),.A(I15598));
INVX1 NOT_2602 (.Y(I9452),.A(g5085));
INVX1 NOT_2603 (.Y(g11182),.A(I16947));
INVX1 NOT_2604 (.Y(g11651),.A(I17755));
INVX1 NOT_2605 (.Y(g7064),.A(I11269));
INVX1 NOT_2606 (.Y(I5210),.A(g58));
INVX1 NOT_2607 (.Y(g2239),.A(I5240));
INVX1 NOT_2608 (.Y(I10180),.A(g6107));
INVX1 NOT_2609 (.Y(g9672),.A(I14805));
INVX1 NOT_2610 (.Y(I13708),.A(g8337));
INVX1 NOT_2611 (.Y(g5774),.A(I9362));
INVX1 NOT_2612 (.Y(g7899),.A(I12683));
INVX1 NOT_2613 (.Y(g3793),.A(g2593));
INVX1 NOT_2614 (.Y(g7464),.A(I11858));
INVX1 NOT_2615 (.Y(I12053),.A(g6928));
INVX1 NOT_2616 (.Y(g8358),.A(I13454));
INVX1 NOT_2617 (.Y(I12809),.A(g7686));
INVX1 NOT_2618 (.Y(g7785),.A(I12520));
INVX1 NOT_2619 (.Y(I16811),.A(g10908));
INVX1 NOT_2620 (.Y(g10551),.A(I16214));
INVX1 NOT_2621 (.Y(I6233),.A(g2299));
INVX1 NOT_2622 (.Y(g2832),.A(I5946));
INVX1 NOT_2623 (.Y(I12466),.A(g7585));
INVX1 NOT_2624 (.Y(g3415),.A(g3121));
INVX1 NOT_2625 (.Y(g3227),.A(I6406));
INVX1 NOT_2626 (.Y(I7825),.A(g3414));
INVX1 NOT_2627 (.Y(g6799),.A(I10807));
INVX1 NOT_2628 (.Y(g2853),.A(g2171));
INVX1 NOT_2629 (.Y(I11043),.A(g6412));
INVX1 NOT_2630 (.Y(I6454),.A(g2368));
INVX1 NOT_2631 (.Y(I13043),.A(g8055));
INVX1 NOT_2632 (.Y(I17216),.A(g11291));
INVX1 NOT_2633 (.Y(g2420),.A(g237));
INVX1 NOT_2634 (.Y(g6674),.A(I10639));
INVX1 NOT_2635 (.Y(I9486),.A(g5066));
INVX1 NOT_2636 (.Y(g11513),.A(I17558));
INVX1 NOT_2637 (.Y(I12177),.A(g7259));
INVX1 NOT_2638 (.Y(g10127),.A(I15383));
INVX1 NOT_2639 (.Y(g3664),.A(g3209));
INVX1 NOT_2640 (.Y(g8275),.A(I13197));
INVX1 NOT_2641 (.Y(g2507),.A(I5584));
INVX1 NOT_2642 (.Y(g8311),.A(I13317));
INVX1 NOT_2643 (.Y(g3246),.A(g2482));
INVX1 NOT_2644 (.Y(I15448),.A(g10056));
INVX1 NOT_2645 (.Y(g5509),.A(g4739));
INVX1 NOT_2646 (.Y(g4326),.A(g3863));
INVX1 NOT_2647 (.Y(I14694),.A(g9259));
INVX1 NOT_2648 (.Y(I7408),.A(g4125));
INVX1 NOT_2649 (.Y(g7237),.A(I11477));
INVX1 NOT_2650 (.Y(g10490),.A(I16105));
INVX1 NOT_2651 (.Y(I9185),.A(g4915));
INVX1 NOT_2652 (.Y(I7336),.A(g3997));
INVX1 NOT_2653 (.Y(g3721),.A(I6891));
INVX1 NOT_2654 (.Y(g11505),.A(I17534));
INVX1 NOT_2655 (.Y(I11602),.A(g6833));
INVX1 NOT_2656 (.Y(I11810),.A(g7246));
INVX1 NOT_2657 (.Y(g11404),.A(I17255));
INVX1 NOT_2658 (.Y(g6132),.A(I9833));
INVX1 NOT_2659 (.Y(g5662),.A(I9147));
INVX1 NOT_2660 (.Y(I6553),.A(g3186));
INVX1 NOT_2661 (.Y(I4850),.A(g1958));
INVX1 NOT_2662 (.Y(g7844),.A(I12631));
INVX1 NOT_2663 (.Y(I17543),.A(g11499));
INVX1 NOT_2664 (.Y(I11068),.A(g6426));
INVX1 NOT_2665 (.Y(I13068),.A(g7906));
INVX1 NOT_2666 (.Y(g6680),.A(I10643));
INVX1 NOT_2667 (.Y(g6209),.A(I9956));
INVX1 NOT_2668 (.Y(g8985),.A(I14376));
INVX1 NOT_2669 (.Y(I11879),.A(g6893));
INVX1 NOT_2670 (.Y(g5994),.A(I9612));
INVX1 NOT_2671 (.Y(g10889),.A(I16629));
INVX1 NOT_2672 (.Y(I16850),.A(g10905));
INVX1 NOT_2673 (.Y(I11970),.A(g6918));
INVX1 NOT_2674 (.Y(g7394),.A(I11778));
INVX1 NOT_2675 (.Y(I10557),.A(g6197));
INVX1 NOT_2676 (.Y(g10354),.A(I15826));
INVX1 NOT_2677 (.Y(g2905),.A(I6068));
INVX1 NOT_2678 (.Y(g7089),.A(I11322));
INVX1 NOT_2679 (.Y(g7731),.A(I12376));
INVX1 NOT_2680 (.Y(g10888),.A(I16626));
INVX1 NOT_2681 (.Y(g6802),.A(I10816));
INVX1 NOT_2682 (.Y(g8239),.A(g7826));
INVX1 NOT_2683 (.Y(g4183),.A(I7366));
INVX1 NOT_2684 (.Y(g9273),.A(I14490));
INVX1 NOT_2685 (.Y(g4608),.A(g3829));
INVX1 NOT_2686 (.Y(g5816),.A(I9424));
INVX1 NOT_2687 (.Y(I5922),.A(g2170));
INVX1 NOT_2688 (.Y(I7465),.A(g3726));
INVX1 NOT_2689 (.Y(g7966),.A(I12762));
INVX1 NOT_2690 (.Y(g2100),.A(I4948));
INVX1 NOT_2691 (.Y(I10278),.A(g5815));
INVX1 NOT_2692 (.Y(g3940),.A(g2920));
INVX1 NOT_2693 (.Y(g6558),.A(I10484));
INVX1 NOT_2694 (.Y(I12009),.A(g6915));
INVX1 NOT_2695 (.Y(I6888),.A(g2960));
INVX1 NOT_2696 (.Y(I8262),.A(g4636));
INVX1 NOT_2697 (.Y(I11967),.A(g6911));
INVX1 NOT_2698 (.Y(g8020),.A(I12862));
INVX1 NOT_2699 (.Y(I10286),.A(g6237));
INVX1 NOT_2700 (.Y(g8420),.A(I13574));
INVX1 NOT_2701 (.Y(I5060),.A(g1191));
INVX1 NOT_2702 (.Y(g10931),.A(g10827));
INVX1 NOT_2703 (.Y(g3388),.A(I6590));
INVX1 NOT_2704 (.Y(I10039),.A(g5718));
INVX1 NOT_2705 (.Y(I14306),.A(g8812));
INVX1 NOT_2706 (.Y(I11459),.A(g6488));
INVX1 NOT_2707 (.Y(g11433),.A(I17350));
INVX1 NOT_2708 (.Y(g9572),.A(I14709));
INVX1 NOT_2709 (.Y(g5685),.A(I9208));
INVX1 NOT_2710 (.Y(g5197),.A(I8611));
INVX1 NOT_2711 (.Y(g5700),.A(I9237));
INVX1 NOT_2712 (.Y(g8794),.A(I14109));
INVX1 NOT_2713 (.Y(g5397),.A(I8835));
INVX1 NOT_2714 (.Y(g2750),.A(I5818));
INVX1 NOT_2715 (.Y(I8889),.A(g4553));
INVX1 NOT_2716 (.Y(g11620),.A(I17678));
INVX1 NOT_2717 (.Y(g10190),.A(I15548));
INVX1 NOT_2718 (.Y(I8476),.A(g4577));
INVX1 NOT_2719 (.Y(g4361),.A(I7648));
INVX1 NOT_2720 (.Y(I9766),.A(g5348));
INVX1 NOT_2721 (.Y(I15811),.A(g10200));
INVX1 NOT_2722 (.Y(g3428),.A(I6639));
INVX1 NOT_2723 (.Y(I7096),.A(g3186));
INVX1 NOT_2724 (.Y(I12454),.A(g7544));
INVX1 NOT_2725 (.Y(I9087),.A(g5113));
INVX1 NOT_2726 (.Y(I9105),.A(g5589));
INVX1 NOT_2727 (.Y(I9305),.A(g4970));
INVX1 NOT_2728 (.Y(I9801),.A(g5416));
INVX1 NOT_2729 (.Y(g3430),.A(I6643));
INVX1 NOT_2730 (.Y(g7814),.A(I12607));
INVX1 NOT_2731 (.Y(I12712),.A(g7441));
INVX1 NOT_2732 (.Y(g11646),.A(I17742));
INVX1 NOT_2733 (.Y(g4051),.A(I7166));
INVX1 NOT_2734 (.Y(I10601),.A(g5996));
INVX1 NOT_2735 (.Y(I13010),.A(g8047));
INVX1 NOT_2736 (.Y(g11343),.A(I17152));
INVX1 NOT_2737 (.Y(I13918),.A(g8451));
INVX1 NOT_2738 (.Y(I16379),.A(g10598));
INVX1 NOT_2739 (.Y(g4127),.A(I7276));
INVX1 NOT_2740 (.Y(g4451),.A(g3638));
INVX1 NOT_2741 (.Y(I15971),.A(g10408));
INVX1 NOT_2742 (.Y(g4327),.A(I7600));
INVX1 NOT_2743 (.Y(I17265),.A(g11352));
INVX1 NOT_2744 (.Y(g7350),.A(I11698));
INVX1 NOT_2745 (.Y(g2040),.A(g1786));
INVX1 NOT_2746 (.Y(g6574),.A(I10514));
INVX1 NOT_2747 (.Y(I12907),.A(g7959));
INVX1 NOT_2748 (.Y(I5995),.A(g2196));
INVX1 NOT_2749 (.Y(I11079),.A(g6649));
INVX1 NOT_2750 (.Y(g10546),.A(I16203));
INVX1 NOT_2751 (.Y(g7038),.A(I11201));
INVX1 NOT_2752 (.Y(I11444),.A(g6653));
INVX1 NOT_2753 (.Y(I17416),.A(g11420));
INVX1 NOT_2754 (.Y(g10211),.A(I15583));
INVX1 NOT_2755 (.Y(g9534),.A(I14687));
INVX1 NOT_2756 (.Y(g9961),.A(I15162));
INVX1 NOT_2757 (.Y(g6714),.A(g5867));
INVX1 NOT_2758 (.Y(g7438),.A(g7232));
INVX1 NOT_2759 (.Y(g7773),.A(I12484));
INVX1 NOT_2760 (.Y(I11599),.A(g6832));
INVX1 NOT_2761 (.Y(g7009),.A(I11152));
INVX1 NOT_2762 (.Y(g11369),.A(I17194));
INVX1 NOT_2763 (.Y(g2123),.A(I5047));
INVX1 NOT_2764 (.Y(I6639),.A(g2632));
INVX1 NOT_2765 (.Y(g4346),.A(I7625));
INVX1 NOT_2766 (.Y(g8515),.A(I13714));
INVX1 NOT_2767 (.Y(g10088),.A(I15317));
INVX1 NOT_2768 (.Y(I8285),.A(g4771));
INVX1 NOT_2769 (.Y(I10937),.A(g6552));
INVX1 NOT_2770 (.Y(I12239),.A(g7073));
INVX1 NOT_2771 (.Y(I5840),.A(g2432));
INVX1 NOT_2772 (.Y(I15368),.A(g9990));
INVX1 NOT_2773 (.Y(I17510),.A(g11481));
INVX1 NOT_2774 (.Y(I16742),.A(g10857));
INVX1 NOT_2775 (.Y(g8100),.A(g7947));
INVX1 NOT_2776 (.Y(I16944),.A(g11079));
INVX1 NOT_2777 (.Y(g3910),.A(g3015));
INVX1 NOT_2778 (.Y(I13086),.A(g7924));
INVX1 NOT_2779 (.Y(g7769),.A(I12472));
INVX1 NOT_2780 (.Y(I15412),.A(g10075));
INVX1 NOT_2781 (.Y(g3638),.A(I6821));
INVX1 NOT_2782 (.Y(I8139),.A(g3681));
INVX1 NOT_2783 (.Y(g7212),.A(I11444));
INVX1 NOT_2784 (.Y(g5723),.A(I9265));
INVX1 NOT_2785 (.Y(I14884),.A(g9454));
INVX1 NOT_2786 (.Y(g11412),.A(I17277));
INVX1 NOT_2787 (.Y(I11817),.A(g7246));
INVX1 NOT_2788 (.Y(I10168),.A(g5982));
INVX1 NOT_2789 (.Y(g5101),.A(I8473));
INVX1 NOT_2790 (.Y(g5817),.A(I9427));
INVX1 NOT_2791 (.Y(I11322),.A(g6652));
INVX1 NOT_2792 (.Y(g7918),.A(g7505));
INVX1 NOT_2793 (.Y(g5301),.A(g4373));
INVX1 NOT_2794 (.Y(g7967),.A(I12765));
INVX1 NOT_2795 (.Y(g6262),.A(I10045));
INVX1 NOT_2796 (.Y(I15229),.A(g9968));
INVX1 NOT_2797 (.Y(g2351),.A(I5427));
INVX1 NOT_2798 (.Y(I11159),.A(g6478));
INVX1 NOT_2799 (.Y(g10700),.A(I16379));
INVX1 NOT_2800 (.Y(g2648),.A(I5765));
INVX1 NOT_2801 (.Y(I9491),.A(g5072));
INVX1 NOT_2802 (.Y(g10126),.A(I15380));
INVX1 NOT_2803 (.Y(I8024),.A(g4117));
INVX1 NOT_2804 (.Y(I11901),.A(g6897));
INVX1 NOT_2805 (.Y(I16802),.A(g10902));
INVX1 NOT_2806 (.Y(g2530),.A(I5641));
INVX1 NOT_2807 (.Y(g6736),.A(I10739));
INVX1 NOT_2808 (.Y(I13125),.A(g7975));
INVX1 NOT_2809 (.Y(g8750),.A(I14045));
INVX1 NOT_2810 (.Y(I10666),.A(g6042));
INVX1 NOT_2811 (.Y(g4508),.A(g3946));
INVX1 NOT_2812 (.Y(g10250),.A(g10136));
INVX1 NOT_2813 (.Y(g2655),.A(g2013));
INVX1 NOT_2814 (.Y(g4944),.A(g4430));
INVX1 NOT_2815 (.Y(g4240),.A(g3664));
INVX1 NOT_2816 (.Y(I11783),.A(g7246));
INVX1 NOT_2817 (.Y(I16793),.A(g11014));
INVX1 NOT_2818 (.Y(I7342),.A(g4011));
INVX1 NOT_2819 (.Y(I9602),.A(g5013));
INVX1 NOT_2820 (.Y(g4472),.A(I7847));
INVX1 NOT_2821 (.Y(I10015),.A(g5641));
INVX1 NOT_2822 (.Y(I5704),.A(g2056));
INVX1 NOT_2823 (.Y(g7993),.A(I12813));
INVX1 NOT_2824 (.Y(I7255),.A(g3227));
INVX1 NOT_2825 (.Y(g6076),.A(I9717));
INVX1 NOT_2826 (.Y(I4906),.A(g119));
INVX1 NOT_2827 (.Y(I11656),.A(g7122));
INVX1 NOT_2828 (.Y(I6049),.A(g2219));
INVX1 NOT_2829 (.Y(g5751),.A(I9323));
INVX1 NOT_2830 (.Y(g3758),.A(I6955));
INVX1 NOT_2831 (.Y(g3066),.A(g2135));
INVX1 NOT_2832 (.Y(I8231),.A(g4170));
INVX1 NOT_2833 (.Y(g4443),.A(g3359));
INVX1 NOT_2834 (.Y(g10296),.A(I15708));
INVX1 NOT_2835 (.Y(g8440),.A(I13618));
INVX1 NOT_2836 (.Y(I11680),.A(g7064));
INVX1 NOT_2837 (.Y(g8969),.A(I14340));
INVX1 NOT_2838 (.Y(I17116),.A(g11229));
INVX1 NOT_2839 (.Y(g2410),.A(g1453));
INVX1 NOT_2840 (.Y(g9679),.A(g9452));
INVX1 NOT_2841 (.Y(I7726),.A(g3378));
INVX1 NOT_2842 (.Y(g6175),.A(g5320));
INVX1 NOT_2843 (.Y(g4116),.A(I7260));
INVX1 NOT_2844 (.Y(I7154),.A(g2617));
INVX1 NOT_2845 (.Y(g8323),.A(I13351));
INVX1 NOT_2846 (.Y(g6871),.A(g6724));
INVX1 NOT_2847 (.Y(g2884),.A(I6040));
INVX1 NOT_2848 (.Y(I7354),.A(g4066));
INVX1 NOT_2849 (.Y(g2839),.A(I5957));
INVX1 NOT_2850 (.Y(g3365),.A(I6553));
INVX1 NOT_2851 (.Y(g3861),.A(I7054));
INVX1 NOT_2852 (.Y(I6498),.A(g2958));
INVX1 NOT_2853 (.Y(I17746),.A(g11643));
INVX1 NOT_2854 (.Y(g3055),.A(g2135));
INVX1 NOT_2855 (.Y(I5053),.A(g1188));
INVX1 NOT_2856 (.Y(I15959),.A(g10402));
INVX1 NOT_2857 (.Y(g6285),.A(I10114));
INVX1 NOT_2858 (.Y(g11627),.A(I17695));
INVX1 NOT_2859 (.Y(g7921),.A(g7463));
INVX1 NOT_2860 (.Y(g10197),.A(I15565));
INVX1 NOT_2861 (.Y(g5673),.A(I9180));
INVX1 NOT_2862 (.Y(g4347),.A(g3880));
INVX1 NOT_2863 (.Y(I8551),.A(g4342));
INVX1 NOT_2864 (.Y(I10084),.A(g5742));
INVX1 NOT_2865 (.Y(g2172),.A(g43));
INVX1 NOT_2866 (.Y(g3333),.A(g2779));
INVX1 NOT_2867 (.Y(I9415),.A(g5047));
INVX1 NOT_2868 (.Y(g11112),.A(I16897));
INVX1 NOT_2869 (.Y(I17237),.A(g11394));
INVX1 NOT_2870 (.Y(g4681),.A(g3546));
INVX1 NOT_2871 (.Y(g10870),.A(I16580));
INVX1 NOT_2872 (.Y(g11050),.A(I16811));
INVX1 NOT_2873 (.Y(I8499),.A(g4330));
INVX1 NOT_2874 (.Y(I12577),.A(g7532));
INVX1 NOT_2875 (.Y(g8151),.A(g8036));
INVX1 NOT_2876 (.Y(g10527),.A(g10462));
INVX1 NOT_2877 (.Y(g3774),.A(I6999));
INVX1 NOT_2878 (.Y(g8351),.A(I13433));
INVX1 NOT_2879 (.Y(I17340),.A(g11366));
INVX1 NOT_2880 (.Y(g4533),.A(I7938));
INVX1 NOT_2881 (.Y(I13017),.A(g7848));
INVX1 NOT_2882 (.Y(I13364),.A(g8221));
INVX1 NOT_2883 (.Y(I15386),.A(g10101));
INVX1 NOT_2884 (.Y(g6184),.A(I9915));
INVX1 NOT_2885 (.Y(g2235),.A(g96));
INVX1 NOT_2886 (.Y(g2343),.A(g1927));
INVX1 NOT_2887 (.Y(I12439),.A(g7663));
INVX1 NOT_2888 (.Y(g5669),.A(I9168));
INVX1 NOT_2889 (.Y(I10531),.A(g6169));
INVX1 NOT_2890 (.Y(I17684),.A(g11609));
INVX1 NOT_2891 (.Y(g6339),.A(I10240));
INVX1 NOT_2892 (.Y(I14179),.A(g8785));
INVX1 NOT_2893 (.Y(g4210),.A(I7447));
INVX1 NOT_2894 (.Y(I14531),.A(g9273));
INVX1 NOT_2895 (.Y(I7112),.A(g3186));
INVX1 NOT_2896 (.Y(I17142),.A(g11301));
INVX1 NOT_2897 (.Y(g11096),.A(I16879));
INVX1 NOT_2898 (.Y(g7620),.A(I12208));
INVX1 NOT_2899 (.Y(g4596),.A(I8007));
INVX1 NOT_2900 (.Y(g3538),.A(I6726));
INVX1 NOT_2901 (.Y(I6019),.A(g2554));
INVX1 NOT_2902 (.Y(g4013),.A(I7157));
INVX1 NOT_2903 (.Y(g6424),.A(g6140));
INVX1 NOT_2904 (.Y(I16626),.A(g10859));
INVX1 NOT_2905 (.Y(I10186),.A(g6110));
INVX1 NOT_2906 (.Y(g6737),.A(g6016));
INVX1 NOT_2907 (.Y(g10867),.A(I16571));
INVX1 NOT_2908 (.Y(g2334),.A(I5388));
INVX1 NOT_2909 (.Y(g10894),.A(I16644));
INVX1 NOT_2910 (.Y(g6809),.A(I10837));
INVX1 NOT_2911 (.Y(I10685),.A(g6054));
INVX1 NOT_2912 (.Y(g5743),.A(I9311));
INVX1 NOT_2913 (.Y(g4413),.A(I7749));
INVX1 NOT_2914 (.Y(g5890),.A(g5361));
INVX1 NOT_2915 (.Y(I11289),.A(g6508));
INVX1 NOT_2916 (.Y(I6052),.A(g2220));
INVX1 NOT_2917 (.Y(g2548),.A(I5667));
INVX1 NOT_2918 (.Y(I14373),.A(g8956));
INVX1 NOT_2919 (.Y(I11309),.A(g6531));
INVX1 NOT_2920 (.Y(I5929),.A(g2225));
INVX1 NOT_2921 (.Y(I13023),.A(g8050));
INVX1 NOT_2922 (.Y(g8884),.A(I14224));
INVX1 NOT_2923 (.Y(I16298),.A(g10553));
INVX1 NOT_2924 (.Y(I13224),.A(g8261));
INVX1 NOT_2925 (.Y(g7788),.A(I12529));
INVX1 NOT_2926 (.Y(g6077),.A(I9720));
INVX1 NOT_2927 (.Y(g11429),.A(I17340));
INVX1 NOT_2928 (.Y(g5011),.A(I8385));
INVX1 NOT_2929 (.Y(I16775),.A(g10889));
INVX1 NOT_2930 (.Y(g3067),.A(I6273));
INVX1 NOT_2931 (.Y(I13571),.A(g8355));
INVX1 NOT_2932 (.Y(g10315),.A(g10243));
INVX1 NOT_2933 (.Y(g5856),.A(g5245));
INVX1 NOT_2934 (.Y(g5734),.A(I9290));
INVX1 NOT_2935 (.Y(g10819),.A(I16525));
INVX1 NOT_2936 (.Y(g11428),.A(I17337));
INVX1 NOT_2937 (.Y(g10910),.A(I16682));
INVX1 NOT_2938 (.Y(g3290),.A(I6461));
INVX1 NOT_2939 (.Y(I17362),.A(g11376));
INVX1 NOT_2940 (.Y(g10202),.A(g10171));
INVX1 NOT_2941 (.Y(I10334),.A(g6003));
INVX1 NOT_2942 (.Y(g10257),.A(g10197));
INVX1 NOT_2943 (.Y(g4317),.A(I7586));
INVX1 NOT_2944 (.Y(g8278),.A(I13206));
INVX1 NOT_2945 (.Y(I4876),.A(g580));
INVX1 NOT_2946 (.Y(g3093),.A(I6299));
INVX1 NOT_2947 (.Y(g1998),.A(g802));
INVX1 NOT_2948 (.Y(g5474),.A(I8889));
INVX1 NOT_2949 (.Y(g10111),.A(I15347));
INVX1 NOT_2950 (.Y(g7192),.A(g6742));
INVX1 NOT_2951 (.Y(g5992),.A(I9608));
INVX1 NOT_2952 (.Y(g7085),.A(I11318));
INVX1 NOT_2953 (.Y(g3256),.A(I6424));
INVX1 NOT_2954 (.Y(I7746),.A(g3763));
INVX1 NOT_2955 (.Y(g6634),.A(I10589));
INVX1 NOT_2956 (.Y(I9188),.A(g4908));
INVX1 NOT_2957 (.Y(I10762),.A(g6127));
INVX1 NOT_2958 (.Y(g8667),.A(I13952));
INVX1 NOT_2959 (.Y(g3816),.A(g3228));
INVX1 NOT_2960 (.Y(g8143),.A(g8029));
INVX1 NOT_2961 (.Y(I13816),.A(g8559));
INVX1 NOT_2962 (.Y(I15548),.A(g10083));
INVX1 NOT_2963 (.Y(I6504),.A(g3214));
INVX1 NOT_2964 (.Y(I9388),.A(g5576));
INVX1 NOT_2965 (.Y(g8235),.A(g7967));
INVX1 NOT_2966 (.Y(g8343),.A(I13409));
INVX1 NOT_2967 (.Y(g6742),.A(g5830));
INVX1 NOT_2968 (.Y(g11548),.A(g11519));
INVX1 NOT_2969 (.Y(g6104),.A(I9769));
INVX1 NOT_2970 (.Y(I14964),.A(g9762));
INVX1 NOT_2971 (.Y(g10590),.A(I16255));
INVX1 NOT_2972 (.Y(I9216),.A(g4935));
INVX1 NOT_2973 (.Y(I6385),.A(g2260));
INVX1 NOT_2974 (.Y(g6304),.A(I10171));
INVX1 NOT_2975 (.Y(I16856),.A(g10909));
INVX1 NOT_2976 (.Y(g8566),.A(I13791));
INVX1 NOT_2977 (.Y(g6499),.A(g5867));
INVX1 NOT_2978 (.Y(I16261),.A(g10556));
INVX1 NOT_2979 (.Y(g2202),.A(g148));
INVX1 NOT_2980 (.Y(g11504),.A(I17531));
INVX1 NOT_2981 (.Y(g8988),.A(I14385));
INVX1 NOT_2982 (.Y(g4775),.A(I8139));
INVX1 NOT_2983 (.Y(I11752),.A(g7032));
INVX1 NOT_2984 (.Y(g8134),.A(I13005));
INVX1 NOT_2985 (.Y(g7941),.A(g7406));
INVX1 NOT_2986 (.Y(I15317),.A(g10025));
INVX1 NOT_2987 (.Y(I6025),.A(g2259));
INVX1 NOT_2988 (.Y(g2908),.A(I6077));
INVX1 NOT_2989 (.Y(g8334),.A(I13382));
INVX1 NOT_2990 (.Y(g9265),.A(g8892));
INVX1 NOT_2991 (.Y(g6926),.A(I11046));
INVX1 NOT_2992 (.Y(g2094),.A(I4924));
INVX1 NOT_2993 (.Y(I12415),.A(g7631));
INVX1 NOT_2994 (.Y(g11317),.A(I17112));
INVX1 NOT_2995 (.Y(g10094),.A(I15329));
INVX1 NOT_2996 (.Y(g3397),.A(g2896));
INVX1 NOT_2997 (.Y(g8548),.A(g8390));
INVX1 NOT_2998 (.Y(g2518),.A(g590));
INVX1 NOT_2999 (.Y(g4060),.A(g3144));
INVX1 NOT_3000 (.Y(g4460),.A(g3820));
INVX1 NOT_3001 (.Y(I9564),.A(g5109));
INVX1 NOT_3002 (.Y(I7468),.A(g3697));
INVX1 NOT_3003 (.Y(g6273),.A(I10078));
INVX1 NOT_3004 (.Y(I8885),.A(g4548));
INVX1 NOT_3005 (.Y(g8804),.A(I14133));
INVX1 NOT_3006 (.Y(I14543),.A(g9311));
INVX1 NOT_3007 (.Y(I8414),.A(g4293));
INVX1 NOT_3008 (.Y(g10150),.A(I15448));
INVX1 NOT_3009 (.Y(g10801),.A(I16507));
INVX1 NOT_3010 (.Y(I9826),.A(g5390));
INVX1 NOT_3011 (.Y(I10117),.A(g6241));
INVX1 NOT_3012 (.Y(g7708),.A(I12339));
INVX1 NOT_3013 (.Y(I13669),.A(g8294));
INVX1 NOT_3014 (.Y(g10735),.A(I16416));
INVX1 NOT_3015 (.Y(g10877),.A(I16601));
INVX1 NOT_3016 (.Y(g11057),.A(g10937));
INVX1 NOT_3017 (.Y(g7520),.A(I11898));
INVX1 NOT_3018 (.Y(g8792),.A(I14105));
INVX1 NOT_3019 (.Y(I17347),.A(g11373));
INVX1 NOT_3020 (.Y(I7677),.A(g3735));
INVX1 NOT_3021 (.Y(I11668),.A(g7043));
INVX1 NOT_3022 (.Y(g6044),.A(I9665));
INVX1 NOT_3023 (.Y(g2593),.A(g1973));
INVX1 NOT_3024 (.Y(g7031),.A(g6413));
INVX1 NOT_3025 (.Y(g4739),.A(g4117));
INVX1 NOT_3026 (.Y(I8903),.A(g4561));
INVX1 NOT_3027 (.Y(g6444),.A(g6158));
INVX1 NOT_3028 (.Y(g11245),.A(g11112));
INVX1 NOT_3029 (.Y(g7431),.A(I11821));
INVX1 NOT_3030 (.Y(I15323),.A(g10019));
INVX1 NOT_3031 (.Y(g6269),.A(I10066));
INVX1 NOT_3032 (.Y(I15299),.A(g9995));
INVX1 NOT_3033 (.Y(g7812),.A(I12601));
INVX1 NOT_3034 (.Y(g11626),.A(I17692));
INVX1 NOT_3035 (.Y(g9770),.A(g9432));
INVX1 NOT_3036 (.Y(g10196),.A(I15562));
INVX1 NOT_3037 (.Y(I11489),.A(g6569));
INVX1 NOT_3038 (.Y(g10695),.A(I16366));
INVX1 NOT_3039 (.Y(g5688),.A(I9213));
INVX1 NOT_3040 (.Y(g11323),.A(I17124));
INVX1 NOT_3041 (.Y(I13489),.A(g8233));
INVX1 NOT_3042 (.Y(g2965),.A(I6196));
INVX1 NOT_3043 (.Y(I6406),.A(g2339));
INVX1 NOT_3044 (.Y(I5475),.A(g1289));
INVX1 NOT_3045 (.Y(I7716),.A(g3751));
INVX1 NOT_3046 (.Y(g6572),.A(g5805));
INVX1 NOT_3047 (.Y(g6862),.A(g6720));
INVX1 NOT_3048 (.Y(g7376),.A(I11756));
INVX1 NOT_3049 (.Y(I5949),.A(g2540));
INVX1 NOT_3050 (.Y(g10526),.A(g10460));
INVX1 NOT_3051 (.Y(g8313),.A(I13323));
INVX1 NOT_3052 (.Y(I12484),.A(g7580));
INVX1 NOT_3053 (.Y(I14242),.A(g8787));
INVX1 NOT_3054 (.Y(I9108),.A(g5593));
INVX1 NOT_3055 (.Y(I15775),.A(g10253));
INVX1 NOT_3056 (.Y(I13424),.A(g8200));
INVX1 NOT_3057 (.Y(g4479),.A(I7858));
INVX1 NOT_3058 (.Y(g9532),.A(I14681));
INVX1 NOT_3059 (.Y(I9308),.A(g5494));
INVX1 NOT_3060 (.Y(g6712),.A(g5984));
INVX1 NOT_3061 (.Y(I8036),.A(g3820));
INVX1 NOT_3062 (.Y(g4294),.A(g3664));
INVX1 NOT_3063 (.Y(I10123),.A(g5676));
INVX1 NOT_3064 (.Y(g6543),.A(g5888));
INVX1 NOT_3065 (.Y(g4840),.A(I8199));
INVX1 NOT_3066 (.Y(I8436),.A(g4462));
INVX1 NOT_3067 (.Y(g9553),.A(I14694));
INVX1 NOT_3068 (.Y(I5292),.A(g76));
INVX1 NOT_3069 (.Y(I9883),.A(g5557));
INVX1 NOT_3070 (.Y(I14123),.A(g8767));
INVX1 NOT_3071 (.Y(g3723),.A(g3071));
INVX1 NOT_3072 (.Y(g7765),.A(I12460));
INVX1 NOT_3073 (.Y(g7286),.A(I11534));
INVX1 NOT_3074 (.Y(g4190),.A(I7387));
INVX1 NOT_3075 (.Y(I5998),.A(g2197));
INVX1 NOT_3076 (.Y(g4390),.A(g3914));
INVX1 NOT_3077 (.Y(I10807),.A(g6396));
INVX1 NOT_3078 (.Y(g10457),.A(I15962));
INVX1 NOT_3079 (.Y(g3817),.A(I7043));
INVX1 NOT_3080 (.Y(g7911),.A(g7664));
INVX1 NOT_3081 (.Y(I5646),.A(g940));
INVX1 NOT_3082 (.Y(I10974),.A(g6563));
INVX1 NOT_3083 (.Y(g8094),.A(g7987));
INVX1 NOT_3084 (.Y(g2050),.A(g1861));
INVX1 NOT_3085 (.Y(g2641),.A(g1987));
INVX1 NOT_3086 (.Y(I8831),.A(g4480));
INVX1 NOT_3087 (.Y(I15232),.A(g9974));
INVX1 NOT_3088 (.Y(I10639),.A(g5830));
INVX1 NOT_3089 (.Y(I17516),.A(g11483));
INVX1 NOT_3090 (.Y(g2450),.A(g1351));
INVX1 NOT_3091 (.Y(I16432),.A(g10702));
INVX1 NOT_3092 (.Y(g4501),.A(g3946));
INVX1 NOT_3093 (.Y(g8518),.A(I13723));
INVX1 NOT_3094 (.Y(g6729),.A(I10724));
INVX1 NOT_3095 (.Y(g6961),.A(I11115));
INVX1 NOT_3096 (.Y(g8567),.A(I13794));
INVX1 NOT_3097 (.Y(I10293),.A(g5863));
INVX1 NOT_3098 (.Y(g4156),.A(I7295));
INVX1 NOT_3099 (.Y(I11713),.A(g7023));
INVX1 NOT_3100 (.Y(g7733),.A(I12380));
INVX1 NOT_3101 (.Y(I5850),.A(g2273));
INVX1 NOT_3102 (.Y(g7270),.A(I11515));
INVX1 NOT_3103 (.Y(g9990),.A(I15190));
INVX1 NOT_3104 (.Y(g6927),.A(I11049));
INVX1 NOT_3105 (.Y(g3751),.A(I6944));
INVX1 NOT_3106 (.Y(I9165),.A(g5037));
INVX1 NOT_3107 (.Y(I16461),.A(g10735));
INVX1 NOT_3108 (.Y(I9571),.A(g5509));
INVX1 NOT_3109 (.Y(I9365),.A(g5392));
INVX1 NOT_3110 (.Y(g7610),.A(I12180));
INVX1 NOT_3111 (.Y(g2179),.A(g89));
INVX1 NOT_3112 (.Y(g4942),.A(I8308));
INVX1 NOT_3113 (.Y(g9029),.A(I14424));
INVX1 NOT_3114 (.Y(g6014),.A(g5309));
INVX1 NOT_3115 (.Y(g7073),.A(I11296));
INVX1 NOT_3116 (.Y(I12799),.A(g7556));
INVX1 NOT_3117 (.Y(g7796),.A(I12553));
INVX1 NOT_3118 (.Y(I12813),.A(g7688));
INVX1 NOT_3119 (.Y(g6885),.A(I10979));
INVX1 NOT_3120 (.Y(g9429),.A(g9082));
INVX1 NOT_3121 (.Y(g22),.A(I4777));
INVX1 NOT_3122 (.Y(g7473),.A(g7148));
INVX1 NOT_3123 (.Y(I10391),.A(g5838));
INVX1 NOT_3124 (.Y(I17209),.A(g11289));
INVX1 NOT_3125 (.Y(g6660),.A(I10623));
INVX1 NOT_3126 (.Y(I11255),.A(g6547));
INVX1 NOT_3127 (.Y(g10256),.A(g10140));
INVX1 NOT_3128 (.Y(I6173),.A(g2125));
INVX1 NOT_3129 (.Y(g11512),.A(I17555));
INVX1 NOT_3130 (.Y(I13255),.A(g8270));
INVX1 NOT_3131 (.Y(I14391),.A(g8928));
INVX1 NOT_3132 (.Y(I16650),.A(g10776));
INVX1 NOT_3133 (.Y(I6373),.A(g2024));
INVX1 NOT_3134 (.Y(I6091),.A(g2270));
INVX1 NOT_3135 (.Y(g5183),.A(g4640));
INVX1 NOT_3136 (.Y(g7124),.A(I11363));
INVX1 NOT_3137 (.Y(g7980),.A(I12786));
INVX1 NOT_3138 (.Y(g7324),.A(I11620));
INVX1 NOT_3139 (.Y(g10280),.A(g10160));
INVX1 NOT_3140 (.Y(g6903),.A(I11005));
INVX1 NOT_3141 (.Y(g2777),.A(g2276));
INVX1 NOT_3142 (.Y(I5919),.A(g2530));
INVX1 NOT_3143 (.Y(I11188),.A(g6513));
INVX1 NOT_3144 (.Y(g7069),.A(I11286));
INVX1 NOT_3145 (.Y(I12805),.A(g7684));
INVX1 NOT_3146 (.Y(I13188),.A(g8171));
INVX1 NOT_3147 (.Y(g5779),.A(I9371));
INVX1 NOT_3148 (.Y(I13678),.A(g8306));
INVX1 NOT_3149 (.Y(I14579),.A(g9272));
INVX1 NOT_3150 (.Y(g4954),.A(g4509));
INVX1 NOT_3151 (.Y(g4250),.A(g3698));
INVX1 NOT_3152 (.Y(g4163),.A(I7308));
INVX1 NOT_3153 (.Y(I5952),.A(g2506));
INVX1 NOT_3154 (.Y(g2882),.A(I6034));
INVX1 NOT_3155 (.Y(g7540),.A(I11956));
INVX1 NOT_3156 (.Y(g8160),.A(I13057));
INVX1 NOT_3157 (.Y(g4363),.A(I7654));
INVX1 NOT_3158 (.Y(I11686),.A(g7039));
INVX1 NOT_3159 (.Y(I16528),.A(g10732));
INVX1 NOT_3160 (.Y(I7577),.A(g4124));
INVX1 NOT_3161 (.Y(I5276),.A(g1411));
INVX1 NOT_3162 (.Y(g8360),.A(I13460));
INVX1 NOT_3163 (.Y(I16843),.A(g10898));
INVX1 NOT_3164 (.Y(I6007),.A(g2199));
INVX1 NOT_3165 (.Y(g5423),.A(g4300));
INVX1 NOT_3166 (.Y(I13460),.A(g8155));
INVX1 NOT_3167 (.Y(I17453),.A(g11451));
INVX1 NOT_3168 (.Y(I11383),.A(g6385));
INVX1 NOT_3169 (.Y(g2271),.A(g877));
INVX1 NOT_3170 (.Y(g7377),.A(I11759));
INVX1 NOT_3171 (.Y(g7206),.A(I11436));
INVX1 NOT_3172 (.Y(g10157),.A(I15467));
INVX1 NOT_3173 (.Y(g11445),.A(I17384));
INVX1 NOT_3174 (.Y(g6036),.A(I9647));
INVX1 NOT_3175 (.Y(I5561),.A(g869));
INVX1 NOT_3176 (.Y(I13030),.A(g8052));
INVX1 NOT_3177 (.Y(g2611),.A(I5734));
INVX1 NOT_3178 (.Y(g4453),.A(I7810));
INVX1 NOT_3179 (.Y(g8450),.A(I13648));
INVX1 NOT_3180 (.Y(g6178),.A(g4977));
INVX1 NOT_3181 (.Y(I6767),.A(g2914));
INVX1 NOT_3182 (.Y(g11499),.A(I17516));
INVX1 NOT_3183 (.Y(I8495),.A(g4325));
INVX1 NOT_3184 (.Y(g3368),.A(g3138));
INVX1 NOT_3185 (.Y(g9745),.A(g9454));
INVX1 NOT_3186 (.Y(I11065),.A(g6750));
INVX1 NOT_3187 (.Y(I6535),.A(g2826));
INVX1 NOT_3188 (.Y(g1987),.A(g762));
INVX1 NOT_3189 (.Y(g9338),.A(I14519));
INVX1 NOT_3190 (.Y(g7287),.A(I11537));
INVX1 NOT_3191 (.Y(g2799),.A(g2276));
INVX1 NOT_3192 (.Y(g11498),.A(I17513));
INVX1 NOT_3193 (.Y(I5986),.A(g2194));
INVX1 NOT_3194 (.Y(g6135),.A(I9842));
INVX1 NOT_3195 (.Y(g5665),.A(I9156));
INVX1 NOT_3196 (.Y(g9109),.A(I14452));
INVX1 NOT_3197 (.Y(g6335),.A(I10228));
INVX1 NOT_3198 (.Y(I15989),.A(g10417));
INVX1 NOT_3199 (.Y(g9309),.A(g8892));
INVX1 NOT_3200 (.Y(g3531),.A(g2971));
INVX1 NOT_3201 (.Y(I8869),.A(g4421));
INVX1 NOT_3202 (.Y(g5127),.A(I8535));
INVX1 NOT_3203 (.Y(g3458),.A(g3144));
INVX1 NOT_3204 (.Y(g6182),.A(g5446));
INVX1 NOT_3205 (.Y(g6288),.A(I10123));
INVX1 NOT_3206 (.Y(I17274),.A(g11389));
INVX1 NOT_3207 (.Y(g6382),.A(I10278));
INVX1 NOT_3208 (.Y(I9662),.A(g5319));
INVX1 NOT_3209 (.Y(g8179),.A(I13086));
INVX1 NOT_3210 (.Y(g7849),.A(I12644));
INVX1 NOT_3211 (.Y(g10876),.A(I16598));
INVX1 NOT_3212 (.Y(g10885),.A(g10809));
INVX1 NOT_3213 (.Y(g11056),.A(g10950));
INVX1 NOT_3214 (.Y(g3743),.A(I6932));
INVX1 NOT_3215 (.Y(g8379),.A(I13485));
INVX1 NOT_3216 (.Y(g4912),.A(I8282));
INVX1 NOT_3217 (.Y(I14116),.A(g8766));
INVX1 NOT_3218 (.Y(g2997),.A(g2135));
INVX1 NOT_3219 (.Y(g11611),.A(I17657));
INVX1 NOT_3220 (.Y(I12400),.A(g7537));
INVX1 NOT_3221 (.Y(g2541),.A(I5658));
INVX1 NOT_3222 (.Y(g11080),.A(I16853));
INVX1 NOT_3223 (.Y(I7426),.A(g3334));
INVX1 NOT_3224 (.Y(I9290),.A(g5052));
INVX1 NOT_3225 (.Y(g5146),.A(g4596));
INVX1 NOT_3226 (.Y(g10854),.A(g10708));
INVX1 NOT_3227 (.Y(g6805),.A(I10825));
INVX1 NOT_3228 (.Y(g5633),.A(g4388));
INVX1 NOT_3229 (.Y(g3505),.A(I6694));
INVX1 NOT_3230 (.Y(g7781),.A(I12508));
INVX1 NOT_3231 (.Y(I5970),.A(g2185));
INVX1 NOT_3232 (.Y(g6749),.A(I10756));
INVX1 NOT_3233 (.Y(I16708),.A(g10822));
INVX1 NOT_3234 (.Y(g2238),.A(I5237));
INVX1 NOT_3235 (.Y(g11432),.A(I17347));
INVX1 NOT_3236 (.Y(I13837),.A(g8488));
INVX1 NOT_3237 (.Y(g3411),.A(I6616));
INVX1 NOT_3238 (.Y(I9093),.A(g5397));
INVX1 NOT_3239 (.Y(g7900),.A(g7712));
INVX1 NOT_3240 (.Y(I16258),.A(g10555));
INVX1 NOT_3241 (.Y(I4948),.A(g586));
INVX1 NOT_3242 (.Y(g2209),.A(g93));
INVX1 NOT_3243 (.Y(g7797),.A(I12556));
INVX1 NOT_3244 (.Y(I9256),.A(g5078));
INVX1 NOT_3245 (.Y(I8265),.A(g4602));
INVX1 NOT_3246 (.Y(I9816),.A(g5576));
INVX1 NOT_3247 (.Y(g5696),.A(I9229));
INVX1 NOT_3248 (.Y(I15461),.A(g10074));
INVX1 NOT_3249 (.Y(g6947),.A(I11085));
INVX1 NOT_3250 (.Y(I7984),.A(g3621));
INVX1 NOT_3251 (.Y(I5224),.A(g61));
INVX1 NOT_3252 (.Y(I7280),.A(g3208));
INVX1 NOT_3253 (.Y(I10237),.A(g6120));
INVX1 NOT_3254 (.Y(g6798),.A(I10804));
INVX1 NOT_3255 (.Y(I8442),.A(g4464));
INVX1 NOT_3256 (.Y(I12538),.A(g7658));
INVX1 NOT_3257 (.Y(g8271),.A(I13185));
INVX1 NOT_3258 (.Y(g2802),.A(g2276));
INVX1 NOT_3259 (.Y(g11342),.A(I17149));
INVX1 NOT_3260 (.Y(I10340),.A(g6205));
INVX1 NOT_3261 (.Y(g1991),.A(g778));
INVX1 NOT_3262 (.Y(I5120),.A(g622));
INVX1 NOT_3263 (.Y(g3474),.A(I6679));
INVX1 NOT_3264 (.Y(g9449),.A(g9094));
INVX1 NOT_3265 (.Y(g6560),.A(g5759));
INVX1 NOT_3266 (.Y(I14340),.A(g8820));
INVX1 NOT_3267 (.Y(g5753),.A(I9329));
INVX1 NOT_3268 (.Y(I8164),.A(g3566));
INVX1 NOT_3269 (.Y(I15736),.A(g10258));
INVX1 NOT_3270 (.Y(g10456),.A(I15959));
INVX1 NOT_3271 (.Y(g5508),.A(I8929));
INVX1 NOT_3272 (.Y(g11199),.A(g11112));
INVX1 NOT_3273 (.Y(I14684),.A(g9124));
INVX1 NOT_3274 (.Y(g11650),.A(I17752));
INVX1 NOT_3275 (.Y(g7144),.A(I11387));
INVX1 NOT_3276 (.Y(I11617),.A(g6839));
INVX1 NOT_3277 (.Y(g7344),.A(I11680));
INVX1 NOT_3278 (.Y(g5072),.A(I8442));
INVX1 NOT_3279 (.Y(I7636),.A(g3330));
INVX1 NOT_3280 (.Y(I13915),.A(g8451));
INVX1 NOT_3281 (.Y(g5472),.A(I8885));
INVX1 NOT_3282 (.Y(g8981),.A(I14364));
INVX1 NOT_3283 (.Y(I9421),.A(g5063));
INVX1 NOT_3284 (.Y(g8674),.A(I13959));
INVX1 NOT_3285 (.Y(I5789),.A(g2162));
INVX1 NOT_3286 (.Y(g5043),.A(g4840));
INVX1 NOT_3287 (.Y(I11201),.A(g6522));
INVX1 NOT_3288 (.Y(g10314),.A(I15744));
INVX1 NOT_3289 (.Y(g7259),.A(I11494));
INVX1 NOT_3290 (.Y(g5443),.A(I8872));
INVX1 NOT_3291 (.Y(g6208),.A(I9953));
INVX1 NOT_3292 (.Y(I7790),.A(g3782));
INVX1 NOT_3293 (.Y(I16879),.A(g10936));
INVX1 NOT_3294 (.Y(g6302),.A(I10165));
INVX1 NOT_3295 (.Y(g10307),.A(I15729));
INVX1 NOT_3296 (.Y(I15365),.A(g10025));
INVX1 NOT_3297 (.Y(I7061),.A(g3050));
INVX1 NOT_3298 (.Y(g6579),.A(g5949));
INVX1 NOT_3299 (.Y(g5116),.A(g4682));
INVX1 NOT_3300 (.Y(g6869),.A(I10949));
INVX1 NOT_3301 (.Y(g7852),.A(g7479));
INVX1 NOT_3302 (.Y(g7923),.A(g7527));
INVX1 NOT_3303 (.Y(I17164),.A(g11320));
INVX1 NOT_3304 (.Y(I7387),.A(g4083));
INVX1 NOT_3305 (.Y(g10596),.A(I16269));
INVX1 NOT_3306 (.Y(I11467),.A(g6488));
INVX1 NOT_3307 (.Y(I11494),.A(g6574));
INVX1 NOT_3308 (.Y(I13595),.A(g8339));
INVX1 NOT_3309 (.Y(g8132),.A(I12999));
INVX1 NOT_3310 (.Y(g6719),.A(I10710));
INVX1 NOT_3311 (.Y(I12235),.A(g7082));
INVX1 NOT_3312 (.Y(g8332),.A(I13376));
INVX1 NOT_3313 (.Y(g10243),.A(I15635));
INVX1 NOT_3314 (.Y(I11623),.A(g6841));
INVX1 NOT_3315 (.Y(I12683),.A(g7387));
INVX1 NOT_3316 (.Y(I6388),.A(g2329));
INVX1 NOT_3317 (.Y(g8680),.A(I13965));
INVX1 NOT_3318 (.Y(g10431),.A(g10328));
INVX1 NOT_3319 (.Y(I11037),.A(g6629));
INVX1 NOT_3320 (.Y(g8353),.A(I13439));
INVX1 NOT_3321 (.Y(I14130),.A(g8769));
INVX1 NOT_3322 (.Y(I10362),.A(g6224));
INVX1 NOT_3323 (.Y(g2864),.A(g2298));
INVX1 NOT_3324 (.Y(I10165),.A(g5948));
INVX1 NOT_3325 (.Y(I13782),.A(g8515));
INVX1 NOT_3326 (.Y(g6917),.A(I11029));
INVX1 NOT_3327 (.Y(g4894),.A(I8247));
INVX1 NOT_3328 (.Y(I6028),.A(g2208));
INVX1 NOT_3329 (.Y(g10269),.A(g10154));
INVX1 NOT_3330 (.Y(g8802),.A(I14127));
INVX1 NOT_3331 (.Y(I6671),.A(g2757));
INVX1 NOT_3332 (.Y(I6428),.A(g2348));
INVX1 NOT_3333 (.Y(g7886),.A(g7479));
INVX1 NOT_3334 (.Y(g4735),.A(g3546));
INVX1 NOT_3335 (.Y(I17327),.A(g11349));
INVX1 NOT_3336 (.Y(g6265),.A(I10054));
INVX1 NOT_3337 (.Y(g3976),.A(I7109));
INVX1 NOT_3338 (.Y(I6247),.A(g2462));
INVX1 NOT_3339 (.Y(g4782),.A(g4089));
INVX1 NOT_3340 (.Y(I11155),.A(g6470));
INVX1 NOT_3341 (.Y(g10156),.A(I15464));
INVX1 NOT_3342 (.Y(I15708),.A(g10241));
INVX1 NOT_3343 (.Y(I17537),.A(g11497));
INVX1 NOT_3344 (.Y(I13418),.A(g8145));
INVX1 NOT_3345 (.Y(I13822),.A(g8488));
INVX1 NOT_3346 (.Y(g5697),.A(I9232));
INVX1 NOT_3347 (.Y(I10006),.A(g5633));
INVX1 NOT_3348 (.Y(g6442),.A(I10362));
INVX1 NOT_3349 (.Y(g9452),.A(I14645));
INVX1 NOT_3350 (.Y(g7314),.A(I11590));
INVX1 NOT_3351 (.Y(g5210),.A(I8631));
INVX1 NOT_3352 (.Y(I17108),.A(g11225));
INVX1 NOT_3353 (.Y(g11471),.A(I17450));
INVX1 NOT_3354 (.Y(I7345),.A(g4050));
INVX1 NOT_3355 (.Y(I16458),.A(g10734));
INVX1 NOT_3356 (.Y(I8429),.A(g4458));
INVX1 NOT_3357 (.Y(I9605),.A(g5620));
INVX1 NOT_3358 (.Y(g4475),.A(I7852));
INVX1 NOT_3359 (.Y(g5596),.A(I9020));
INVX1 NOT_3360 (.Y(g6164),.A(g5426));
INVX1 NOT_3361 (.Y(I7763),.A(g3769));
INVX1 NOT_3362 (.Y(I7191),.A(g2646));
INVX1 NOT_3363 (.Y(g10734),.A(I16413));
INVX1 NOT_3364 (.Y(I10437),.A(g5755));
INVX1 NOT_3365 (.Y(g10335),.A(I15787));
INVX1 NOT_3366 (.Y(g7650),.A(I12261));
INVX1 NOT_3367 (.Y(g3326),.A(I6495));
INVX1 NOT_3368 (.Y(I15244),.A(g10031));
INVX1 NOT_3369 (.Y(g4292),.A(g3863));
INVX1 NOT_3370 (.Y(g10930),.A(g10827));
INVX1 NOT_3371 (.Y(g11043),.A(I16790));
INVX1 NOT_3372 (.Y(g6454),.A(I10388));
INVX1 NOT_3373 (.Y(g11244),.A(g11112));
INVX1 NOT_3374 (.Y(g4526),.A(I7931));
INVX1 NOT_3375 (.Y(I5478),.A(g1212));
INVX1 NOT_3376 (.Y(g6296),.A(I10147));
INVX1 NOT_3377 (.Y(I11194),.A(g6515));
INVX1 NOT_3378 (.Y(g3760),.A(g3003));
INVX1 NOT_3379 (.Y(g7008),.A(I11149));
INVX1 NOT_3380 (.Y(I13194),.A(g8140));
INVX1 NOT_3381 (.Y(I13589),.A(g8361));
INVX1 NOT_3382 (.Y(g2623),.A(g1999));
INVX1 NOT_3383 (.Y(I17381),.A(g11436));
INVX1 NOT_3384 (.Y(I7536),.A(g4098));
INVX1 NOT_3385 (.Y(I9585),.A(g5241));
INVX1 NOT_3386 (.Y(g2076),.A(I4886));
INVX1 NOT_3387 (.Y(g10131),.A(I15395));
INVX1 NOT_3388 (.Y(g2889),.A(I6049));
INVX1 NOT_3389 (.Y(I11524),.A(g6593));
INVX1 NOT_3390 (.Y(I16598),.A(g10804));
INVX1 NOT_3391 (.Y(g11069),.A(g10974));
INVX1 NOT_3392 (.Y(g4084),.A(g3119));
INVX1 NOT_3393 (.Y(I11836),.A(g7220));
INVX1 NOT_3394 (.Y(I5435),.A(g18));
INVX1 NOT_3395 (.Y(g4603),.A(g3829));
INVX1 NOT_3396 (.Y(g5936),.A(I9564));
INVX1 NOT_3397 (.Y(g7336),.A(I11656));
INVX1 NOT_3398 (.Y(g8600),.A(g8475));
INVX1 NOT_3399 (.Y(I15068),.A(g9710));
INVX1 NOT_3400 (.Y(g7768),.A(I12469));
INVX1 NOT_3401 (.Y(g4439),.A(I7793));
INVX1 NOT_3402 (.Y(g11657),.A(I17773));
INVX1 NOT_3403 (.Y(g5117),.A(g4682));
INVX1 NOT_3404 (.Y(g6553),.A(I10477));
INVX1 NOT_3405 (.Y(g8714),.A(I14005));
INVX1 NOT_3406 (.Y(g11068),.A(g10974));
INVX1 NOT_3407 (.Y(I7858),.A(g3631));
INVX1 NOT_3408 (.Y(I11477),.A(g6488));
INVX1 NOT_3409 (.Y(g7594),.A(I12120));
INVX1 NOT_3410 (.Y(g10487),.A(I16098));
INVX1 NOT_3411 (.Y(g7972),.A(I12770));
INVX1 NOT_3412 (.Y(g2175),.A(g44));
INVX1 NOT_3413 (.Y(I11119),.A(g6461));
INVX1 NOT_3414 (.Y(g9025),.A(I14412));
INVX1 NOT_3415 (.Y(g2871),.A(I6013));
INVX1 NOT_3416 (.Y(g10619),.A(I16292));
INVX1 NOT_3417 (.Y(I12759),.A(g7702));
INVX1 NOT_3418 (.Y(I7757),.A(g3767));
INVX1 NOT_3419 (.Y(I16817),.A(g10912));
INVX1 NOT_3420 (.Y(I9673),.A(g5182));
INVX1 NOT_3421 (.Y(I14236),.A(g8802));
INVX1 NOT_3422 (.Y(g7806),.A(I12583));
INVX1 NOT_3423 (.Y(I10952),.A(g6556));
INVX1 NOT_3424 (.Y(g3220),.A(I6398));
INVX1 NOT_3425 (.Y(I8109),.A(g3622));
INVX1 NOT_3426 (.Y(g2651),.A(g2007));
INVX1 NOT_3427 (.Y(I6217),.A(g2302));
INVX1 NOT_3428 (.Y(g4583),.A(g3880));
INVX1 NOT_3429 (.Y(g6412),.A(I10322));
INVX1 NOT_3430 (.Y(I17390),.A(g11430));
INVX1 NOT_3431 (.Y(g10279),.A(g10158));
INVX1 NOT_3432 (.Y(g7065),.A(I11272));
INVX1 NOT_3433 (.Y(I7315),.A(g2891));
INVX1 NOT_3434 (.Y(g6389),.A(I10289));
INVX1 NOT_3435 (.Y(I7642),.A(g3440));
INVX1 NOT_3436 (.Y(I9168),.A(g5040));
INVX1 NOT_3437 (.Y(g6706),.A(I10685));
INVX1 NOT_3438 (.Y(I9669),.A(g5426));
INVX1 NOT_3439 (.Y(g7887),.A(g7693));
INVX1 NOT_3440 (.Y(g7122),.A(I11357));
INVX1 NOT_3441 (.Y(I15792),.A(g10279));
INVX1 NOT_3442 (.Y(I9368),.A(g5288));
INVX1 NOT_3443 (.Y(g7322),.A(I11614));
INVX1 NOT_3444 (.Y(g4919),.A(I8290));
INVX1 NOT_3445 (.Y(I10063),.A(g5766));
INVX1 NOT_3446 (.Y(g6990),.A(I11132));
INVX1 NOT_3447 (.Y(I7447),.A(g3694));
INVX1 NOT_3448 (.Y(g10278),.A(g10182));
INVX1 NOT_3449 (.Y(g3977),.A(I7112));
INVX1 NOT_3450 (.Y(I6861),.A(g2942));
INVX1 NOT_3451 (.Y(g6888),.A(I10984));
INVX1 NOT_3452 (.Y(I16656),.A(g10791));
INVX1 NOT_3453 (.Y(I9531),.A(g5004));
INVX1 NOT_3454 (.Y(g6171),.A(g5446));
INVX1 NOT_3455 (.Y(g2184),.A(g1806));
INVX1 NOT_3456 (.Y(I16295),.A(g10552));
INVX1 NOT_3457 (.Y(I9458),.A(g5091));
INVX1 NOT_3458 (.Y(g3161),.A(I6367));
INVX1 NOT_3459 (.Y(I11704),.A(g7008));
INVX1 NOT_3460 (.Y(I12849),.A(g7632));
INVX1 NOT_3461 (.Y(I6055),.A(g2569));
INVX1 NOT_3462 (.Y(I17522),.A(g11485));
INVX1 NOT_3463 (.Y(g2339),.A(I5399));
INVX1 NOT_3464 (.Y(g7033),.A(I11188));
INVX1 NOT_3465 (.Y(g10039),.A(I15244));
INVX1 NOT_3466 (.Y(I10873),.A(g6331));
INVX1 NOT_3467 (.Y(g6956),.A(I11106));
INVX1 NOT_3468 (.Y(g5597),.A(I9023));
INVX1 NOT_3469 (.Y(I14873),.A(g9525));
INVX1 NOT_3470 (.Y(I7654),.A(g3728));
INVX1 NOT_3471 (.Y(I13809),.A(g8480));
INVX1 NOT_3472 (.Y(I6133),.A(g2253));
INVX1 NOT_3473 (.Y(g3051),.A(g2135));
INVX1 NOT_3474 (.Y(g2838),.A(g2165));
INVX1 NOT_3475 (.Y(g8076),.A(I12930));
INVX1 NOT_3476 (.Y(g2024),.A(g1718));
INVX1 NOT_3477 (.Y(I15458),.A(g10069));
INVX1 NOT_3478 (.Y(I13466),.A(g8160));
INVX1 NOT_3479 (.Y(I9505),.A(g5088));
INVX1 NOT_3480 (.Y(g6281),.A(I10102));
INVX1 NOT_3481 (.Y(g8476),.A(I13674));
INVX1 NOT_3482 (.Y(g3327),.A(I6498));
INVX1 NOT_3483 (.Y(g2424),.A(g1690));
INVX1 NOT_3484 (.Y(I8449),.A(g4469));
INVX1 NOT_3485 (.Y(I12652),.A(g7458));
INVX1 NOT_3486 (.Y(g9766),.A(g9432));
INVX1 NOT_3487 (.Y(g2809),.A(I5909));
INVX1 NOT_3488 (.Y(g5784),.A(I9380));
INVX1 NOT_3489 (.Y(g4004),.A(I7140));
INVX1 NOT_3490 (.Y(I9734),.A(g5257));
INVX1 NOT_3491 (.Y(I13036),.A(g8053));
INVX1 NOT_3492 (.Y(I5002),.A(g1173));
INVX1 NOT_3493 (.Y(I8865),.A(g4518));
INVX1 NOT_3494 (.Y(g7550),.A(g6974));
INVX1 NOT_3495 (.Y(g6297),.A(I10150));
INVX1 NOT_3496 (.Y(I11560),.A(g7037));
INVX1 NOT_3497 (.Y(g10187),.A(I15539));
INVX1 NOT_3498 (.Y(I6196),.A(g2462));
INVX1 NOT_3499 (.Y(I5824),.A(g2502));
INVX1 NOT_3500 (.Y(g7845),.A(I12634));
INVX1 NOT_3501 (.Y(I10834),.A(g6715));
INVX1 NOT_3502 (.Y(g8871),.A(I14185));
INVX1 NOT_3503 (.Y(g8375),.A(I13475));
INVX1 NOT_3504 (.Y(I15545),.A(g10075));
INVX1 NOT_3505 (.Y(g3633),.A(I6802));
INVX1 NOT_3506 (.Y(I15079),.A(g9745));
INVX1 NOT_3507 (.Y(I8098),.A(g3583));
INVX1 NOT_3508 (.Y(g2077),.A(g219));
INVX1 NOT_3509 (.Y(g2231),.A(I5218));
INVX1 NOT_3510 (.Y(g7195),.A(I11417));
INVX1 NOT_3511 (.Y(g11545),.A(g11519));
INVX1 NOT_3512 (.Y(g11079),.A(I16850));
INVX1 NOT_3513 (.Y(g11444),.A(I17381));
INVX1 NOT_3514 (.Y(g5937),.A(I9567));
INVX1 NOT_3515 (.Y(g7395),.A(g6941));
INVX1 NOT_3516 (.Y(I13642),.A(g8378));
INVX1 NOT_3517 (.Y(g7337),.A(I11659));
INVX1 NOT_3518 (.Y(g3103),.A(g2391));
INVX1 NOT_3519 (.Y(I9074),.A(g4764));
INVX1 NOT_3520 (.Y(g7913),.A(g7467));
INVX1 NOT_3521 (.Y(I6538),.A(g2827));
INVX1 NOT_3522 (.Y(g2523),.A(I5632));
INVX1 NOT_3523 (.Y(I7272),.A(g3253));
INVX1 NOT_3524 (.Y(g2643),.A(g1989));
INVX1 NOT_3525 (.Y(I9992),.A(g5633));
INVX1 NOT_3526 (.Y(g10143),.A(I15427));
INVX1 NOT_3527 (.Y(g5668),.A(I9165));
INVX1 NOT_3528 (.Y(g11078),.A(I16847));
INVX1 NOT_3529 (.Y(g6338),.A(I10237));
INVX1 NOT_3530 (.Y(I15598),.A(g10170));
INVX1 NOT_3531 (.Y(I10021),.A(g5692));
INVX1 NOT_3532 (.Y(g5840),.A(g5320));
INVX1 NOT_3533 (.Y(g4970),.A(g4411));
INVX1 NOT_3534 (.Y(g8500),.A(I13695));
INVX1 NOT_3535 (.Y(I7612),.A(g3817));
INVX1 NOT_3536 (.Y(g11598),.A(I17642));
INVX1 NOT_3537 (.Y(I7017),.A(g3068));
INVX1 NOT_3538 (.Y(g6109),.A(g5052));
INVX1 NOT_3539 (.Y(I12406),.A(g7464));
INVX1 NOT_3540 (.Y(g6309),.A(I10186));
INVX1 NOT_3541 (.Y(g11086),.A(I16867));
INVX1 NOT_3542 (.Y(g7807),.A(I12586));
INVX1 NOT_3543 (.Y(I7417),.A(g4160));
INVX1 NOT_3544 (.Y(g3732),.A(I6914));
INVX1 NOT_3545 (.Y(I17252),.A(g11343));
INVX1 NOT_3546 (.Y(g10169),.A(I15503));
INVX1 NOT_3547 (.Y(I7935),.A(g3440));
INVX1 NOT_3548 (.Y(I9080),.A(g4775));
INVX1 NOT_3549 (.Y(g8184),.A(I13105));
INVX1 NOT_3550 (.Y(g10884),.A(g10809));
INVX1 NOT_3551 (.Y(g6808),.A(I10834));
INVX1 NOT_3552 (.Y(I15817),.A(g10199));
INVX1 NOT_3553 (.Y(I9863),.A(g5557));
INVX1 NOT_3554 (.Y(g8139),.A(g8025));
INVX1 NOT_3555 (.Y(I16289),.A(g10541));
INVX1 NOT_3556 (.Y(g8339),.A(I13397));
INVX1 NOT_3557 (.Y(g2742),.A(I5798));
INVX1 NOT_3558 (.Y(g3944),.A(g2920));
INVX1 NOT_3559 (.Y(g10168),.A(I15500));
INVX1 NOT_3560 (.Y(I10607),.A(g5763));
INVX1 NOT_3561 (.Y(g6707),.A(g5949));
INVX1 NOT_3562 (.Y(I13630),.A(g8334));
INVX1 NOT_3563 (.Y(g2304),.A(I5348));
INVX1 NOT_3564 (.Y(g11322),.A(I17121));
INVX1 NOT_3565 (.Y(g9091),.A(g8892));
INVX1 NOT_3566 (.Y(g4320),.A(g4013));
INVX1 NOT_3567 (.Y(I15977),.A(g10411));
INVX1 NOT_3568 (.Y(g11159),.A(g10950));
INVX1 NOT_3569 (.Y(I10274),.A(g5811));
INVX1 NOT_3570 (.Y(I11166),.A(g6480));
INVX1 NOT_3571 (.Y(I11665),.A(g7038));
INVX1 NOT_3572 (.Y(I16571),.A(g10819));
INVX1 NOT_3573 (.Y(I13166),.A(g8009));
INVX1 NOT_3574 (.Y(I7330),.A(g3761));
INVX1 NOT_3575 (.Y(I8268),.A(g4674));
INVX1 NOT_3576 (.Y(g8424),.A(I13586));
INVX1 NOT_3577 (.Y(I5064),.A(g1690));
INVX1 NOT_3578 (.Y(g8795),.A(I14112));
INVX1 NOT_3579 (.Y(g10217),.A(I15589));
INVX1 NOT_3580 (.Y(g7142),.A(I11383));
INVX1 NOT_3581 (.Y(I6256),.A(g2462));
INVX1 NOT_3582 (.Y(g4277),.A(g3688));
INVX1 NOT_3583 (.Y(g6201),.A(I9938));
INVX1 NOT_3584 (.Y(g7342),.A(I11674));
INVX1 NOT_3585 (.Y(I11008),.A(g6795));
INVX1 NOT_3586 (.Y(g6957),.A(I11109));
INVX1 NOT_3587 (.Y(I15353),.A(g10007));
INVX1 NOT_3588 (.Y(g2754),.A(I5830));
INVX1 NOT_3589 (.Y(g4906),.A(I8275));
INVX1 NOT_3590 (.Y(g7815),.A(I12610));
INVX1 NOT_3591 (.Y(g11656),.A(I17770));
INVX1 NOT_3592 (.Y(g4789),.A(g3337));
INVX1 NOT_3593 (.Y(I7800),.A(g3791));
INVX1 NOT_3594 (.Y(g10486),.A(I16095));
INVX1 NOT_3595 (.Y(g11353),.A(I17176));
INVX1 NOT_3596 (.Y(g8077),.A(I12933));
INVX1 NOT_3597 (.Y(I15823),.A(g10201));
INVX1 NOT_3598 (.Y(g6449),.A(g6172));
INVX1 NOT_3599 (.Y(I13485),.A(g8194));
INVX1 NOT_3600 (.Y(g2273),.A(g881));
INVX1 NOT_3601 (.Y(g8477),.A(g8317));
INVX1 NOT_3602 (.Y(g6575),.A(g5949));
INVX1 NOT_3603 (.Y(g7692),.A(g7148));
INVX1 NOT_3604 (.Y(I12613),.A(g7525));
INVX1 NOT_3605 (.Y(g8523),.A(I13732));
INVX1 NOT_3606 (.Y(I6381),.A(g2257));
INVX1 NOT_3607 (.Y(g9767),.A(I14914));
INVX1 NOT_3608 (.Y(g7097),.A(I11330));
INVX1 NOT_3609 (.Y(I9688),.A(g5201));
INVX1 NOT_3610 (.Y(g7726),.A(I12363));
INVX1 NOT_3611 (.Y(I9857),.A(g5269));
INVX1 NOT_3612 (.Y(I13454),.A(g8183));
INVX1 NOT_3613 (.Y(g2613),.A(I5740));
INVX1 NOT_3614 (.Y(g7497),.A(g7148));
INVX1 NOT_3615 (.Y(g9535),.A(I14690));
INVX1 NOT_3616 (.Y(g6715),.A(I10702));
INVX1 NOT_3617 (.Y(g2044),.A(I4850));
INVX1 NOT_3618 (.Y(g7354),.A(I11710));
INVX1 NOT_3619 (.Y(g10580),.A(g10530));
INVX1 NOT_3620 (.Y(I10153),.A(g5947));
INVX1 NOT_3621 (.Y(g2444),.A(g876));
INVX1 NOT_3622 (.Y(I5237),.A(g1107));
INVX1 NOT_3623 (.Y(g5032),.A(I8403));
INVX1 NOT_3624 (.Y(g2269),.A(I5308));
INVX1 NOT_3625 (.Y(g10223),.A(I15595));
INVX1 NOT_3626 (.Y(I7213),.A(g2635));
INVX1 NOT_3627 (.Y(g9261),.A(g8892));
INVX1 NOT_3628 (.Y(I6421),.A(g2346));
INVX1 NOT_3629 (.Y(g4299),.A(g4144));
INVX1 NOT_3630 (.Y(I14409),.A(g8938));
INVX1 NOT_3631 (.Y(I12463),.A(g7579));
INVX1 NOT_3632 (.Y(g3697),.A(I6856));
INVX1 NOT_3633 (.Y(g8099),.A(g7990));
INVX1 NOT_3634 (.Y(I8385),.A(g4238));
INVX1 NOT_3635 (.Y(I14136),.A(g8775));
INVX1 NOT_3636 (.Y(g8304),.A(I13280));
INVX1 NOT_3637 (.Y(g3914),.A(g3015));
INVX1 NOT_3638 (.Y(I9126),.A(g4891));
INVX1 NOT_3639 (.Y(I13239),.A(g8266));
INVX1 NOT_3640 (.Y(g10110),.A(I15344));
INVX1 NOT_3641 (.Y(g11631),.A(I17707));
INVX1 NOT_3642 (.Y(I9326),.A(g5320));
INVX1 NOT_3643 (.Y(g2543),.A(I5662));
INVX1 NOT_3644 (.Y(g6584),.A(I10538));
INVX1 NOT_3645 (.Y(g11017),.A(I16742));
INVX1 NOT_3646 (.Y(g6539),.A(I10461));
INVX1 NOT_3647 (.Y(g6896),.A(I10996));
INVX1 NOT_3648 (.Y(g5568),.A(I8985));
INVX1 NOT_3649 (.Y(g10321),.A(I15759));
INVX1 NOT_3650 (.Y(I5089),.A(g1854));
INVX1 NOT_3651 (.Y(I5731),.A(g2089));
INVX1 NOT_3652 (.Y(I11238),.A(g6543));
INVX1 NOT_3653 (.Y(I17213),.A(g11290));
INVX1 NOT_3654 (.Y(g7783),.A(I12514));
INVX1 NOT_3655 (.Y(g10179),.A(g10041));
INVX1 NOT_3656 (.Y(g10531),.A(g10471));
INVX1 NOT_3657 (.Y(g7979),.A(I12783));
INVX1 NOT_3658 (.Y(g3413),.A(g2896));
INVX1 NOT_3659 (.Y(g5912),.A(I9544));
INVX1 NOT_3660 (.Y(g7312),.A(I11584));
INVX1 NOT_3661 (.Y(I7166),.A(g2620));
INVX1 NOT_3662 (.Y(I5966),.A(g2541));
INVX1 NOT_3663 (.Y(g10178),.A(I15526));
INVX1 NOT_3664 (.Y(I7366),.A(g4012));
INVX1 NOT_3665 (.Y(g4738),.A(g3440));
INVX1 NOT_3666 (.Y(I13941),.A(g8488));
INVX1 NOT_3667 (.Y(I13382),.A(g8134));
INVX1 NOT_3668 (.Y(g6268),.A(I10063));
INVX1 NOT_3669 (.Y(I11519),.A(g6591));
INVX1 NOT_3670 (.Y(I11176),.A(g6501));
INVX1 NOT_3671 (.Y(g10186),.A(I15536));
INVX1 NOT_3672 (.Y(g7001),.A(I11140));
INVX1 NOT_3673 (.Y(g8273),.A(I13191));
INVX1 NOT_3674 (.Y(g10676),.A(g10570));
INVX1 NOT_3675 (.Y(g6419),.A(I10331));
INVX1 NOT_3676 (.Y(I10891),.A(g6334));
INVX1 NOT_3677 (.Y(I13185),.A(g8192));
INVX1 NOT_3678 (.Y(g11289),.A(I17070));
INVX1 NOT_3679 (.Y(I7456),.A(g3716));
INVX1 NOT_3680 (.Y(g1993),.A(g786));
INVX1 NOT_3681 (.Y(g3820),.A(I7048));
INVX1 NOT_3682 (.Y(g7676),.A(I12303));
INVX1 NOT_3683 (.Y(g4140),.A(I7284));
INVX1 NOT_3684 (.Y(g6052),.A(g5426));
INVX1 NOT_3685 (.Y(g11309),.A(I17096));
INVX1 NOT_3686 (.Y(g4078),.A(I7205));
INVX1 NOT_3687 (.Y(I12514),.A(g7735));
INVX1 NOT_3688 (.Y(g8613),.A(g8484));
INVX1 NOT_3689 (.Y(I16525),.A(g10719));
INVX1 NOT_3690 (.Y(I7348),.A(g4056));
INVX1 NOT_3691 (.Y(g6452),.A(I10384));
INVX1 NOT_3692 (.Y(I9383),.A(g5296));
INVX1 NOT_3693 (.Y(I9608),.A(g5127));
INVX1 NOT_3694 (.Y(I15308),.A(g10019));
INVX1 NOT_3695 (.Y(g7329),.A(I11635));
INVX1 NOT_3696 (.Y(g4478),.A(g3820));
INVX1 NOT_3697 (.Y(g7761),.A(I12448));
INVX1 NOT_3698 (.Y(g2014),.A(g1104));
INVX1 NOT_3699 (.Y(g4907),.A(I8278));
INVX1 NOT_3700 (.Y(g8444),.A(I13630));
INVX1 NOT_3701 (.Y(g2885),.A(I6043));
INVX1 NOT_3702 (.Y(I9779),.A(g5391));
INVX1 NOT_3703 (.Y(g2946),.A(I6133));
INVX1 NOT_3704 (.Y(g4435),.A(g3914));
INVX1 NOT_3705 (.Y(I9023),.A(g4727));
INVX1 NOT_3706 (.Y(g8983),.A(I14370));
INVX1 NOT_3707 (.Y(g4082),.A(I7213));
INVX1 NOT_3708 (.Y(I12421),.A(g7634));
INVX1 NOT_3709 (.Y(I8406),.A(g4274));
INVX1 NOT_3710 (.Y(I5254),.A(g1700));
INVX1 NOT_3711 (.Y(I14109),.A(g8765));
INVX1 NOT_3712 (.Y(g8572),.A(I13809));
INVX1 NOT_3713 (.Y(g7727),.A(I12366));
INVX1 NOT_3714 (.Y(I7964),.A(g3433));
INVX1 NOT_3715 (.Y(g2903),.A(g2166));
INVX1 NOT_3716 (.Y(I7260),.A(g2844));
INVX1 NOT_3717 (.Y(I14537),.A(g9308));
INVX1 NOT_3718 (.Y(I10108),.A(g5743));
INVX1 NOT_3719 (.Y(g6086),.A(I9737));
INVX1 NOT_3720 (.Y(g8712),.A(g8680));
INVX1 NOT_3721 (.Y(g11495),.A(I17500));
INVX1 NOT_3722 (.Y(I12012),.A(g6916));
INVX1 NOT_3723 (.Y(I9588),.A(g5114));
INVX1 NOT_3724 (.Y(g7746),.A(I12403));
INVX1 NOT_3725 (.Y(I8487),.A(g4526));
INVX1 NOT_3726 (.Y(I5438),.A(g18));
INVX1 NOT_3727 (.Y(g3775),.A(I7002));
INVX1 NOT_3728 (.Y(g7221),.A(I11459));
INVX1 NOT_3729 (.Y(I17350),.A(g11377));
INVX1 NOT_3730 (.Y(I14303),.A(g8811));
INVX1 NOT_3731 (.Y(g6385),.A(g6119));
INVX1 NOT_3732 (.Y(g6881),.A(I10971));
INVX1 NOT_3733 (.Y(I12541),.A(g7662));
INVX1 NOT_3734 (.Y(g7703),.A(g7085));
INVX1 NOT_3735 (.Y(I9665),.A(g5174));
INVX1 NOT_3736 (.Y(I15752),.A(g10264));
INVX1 NOT_3737 (.Y(g4915),.A(g4413));
INVX1 NOT_3738 (.Y(g2178),.A(g45));
INVX1 NOT_3739 (.Y(g2436),.A(I5525));
INVX1 NOT_3740 (.Y(I15374),.A(g10007));
INVX1 NOT_3741 (.Y(g9028),.A(I14421));
INVX1 NOT_3742 (.Y(g8729),.A(g8595));
INVX1 NOT_3743 (.Y(g8961),.A(I14330));
INVX1 NOT_3744 (.Y(I4900),.A(g583));
INVX1 NOT_3745 (.Y(I11501),.A(g6581));
INVX1 NOT_3746 (.Y(I16610),.A(g10792));
INVX1 NOT_3747 (.Y(g9671),.A(I14802));
INVX1 NOT_3748 (.Y(I17152),.A(g11308));
INVX1 NOT_3749 (.Y(g3060),.A(g2135));
INVX1 NOT_3750 (.Y(I13729),.A(g8290));
INVX1 NOT_3751 (.Y(I13577),.A(g8330));
INVX1 NOT_3752 (.Y(I10381),.A(g5847));
INVX1 NOT_3753 (.Y(g4214),.A(I7459));
INVX1 NOT_3754 (.Y(I16255),.A(g10554));
INVX1 NOT_3755 (.Y(I14982),.A(g9672));
INVX1 NOT_3756 (.Y(g6425),.A(g6141));
INVX1 NOT_3757 (.Y(I11728),.A(g7010));
INVX1 NOT_3758 (.Y(g11643),.A(I17733));
INVX1 NOT_3759 (.Y(g2135),.A(I5064));
INVX1 NOT_3760 (.Y(I16679),.A(g10784));
INVX1 NOT_3761 (.Y(g2335),.A(I5391));
INVX1 NOT_3762 (.Y(g5683),.A(I9202));
INVX1 NOT_3763 (.Y(I13439),.A(g8187));
INVX1 NOT_3764 (.Y(I9346),.A(g5281));
INVX1 NOT_3765 (.Y(I7118),.A(g2979));
INVX1 NOT_3766 (.Y(g4310),.A(I7577));
INVX1 NOT_3767 (.Y(g2382),.A(g599));
INVX1 NOT_3768 (.Y(I7318),.A(g3266));
INVX1 NOT_3769 (.Y(I12829),.A(g7680));
INVX1 NOT_3770 (.Y(I16124),.A(g10396));
INVX1 NOT_3771 (.Y(g10909),.A(I16679));
INVX1 NOT_3772 (.Y(I12535),.A(g7656));
INVX1 NOT_3773 (.Y(g5778),.A(I9368));
INVX1 NOT_3774 (.Y(I10174),.A(g5994));
INVX1 NOT_3775 (.Y(I15669),.A(g10194));
INVX1 NOT_3776 (.Y(g10543),.A(I16196));
INVX1 NOT_3777 (.Y(g3784),.A(g2586));
INVX1 NOT_3778 (.Y(I17413),.A(g11425));
INVX1 NOT_3779 (.Y(g5894),.A(g5361));
INVX1 NOT_3780 (.Y(g9826),.A(I14979));
INVX1 NOT_3781 (.Y(g10117),.A(I15359));
INVX1 NOT_3782 (.Y(g8660),.A(I13945));
INVX1 NOT_3783 (.Y(g8946),.A(I14295));
INVX1 NOT_3784 (.Y(g10908),.A(I16676));
INVX1 NOT_3785 (.Y(g2916),.A(I6097));
INVX1 NOT_3786 (.Y(I7843),.A(g3440));
INVX1 NOT_3787 (.Y(g2022),.A(g1346));
INVX1 NOT_3788 (.Y(g5735),.A(I9293));
INVX1 NOT_3789 (.Y(I15392),.A(g10104));
INVX1 NOT_3790 (.Y(g7677),.A(g7148));
INVX1 NOT_3791 (.Y(g2749),.A(I5815));
INVX1 NOT_3792 (.Y(g3995),.A(g3121));
INVX1 NOT_3793 (.Y(g3937),.A(I7086));
INVX1 NOT_3794 (.Y(I10840),.A(g6719));
INVX1 NOT_3795 (.Y(g9741),.A(I14888));
INVX1 NOT_3796 (.Y(g4002),.A(g3121));
INVX1 NOT_3797 (.Y(I7393),.A(g4096));
INVX1 NOT_3798 (.Y(I16938),.A(g11086));
INVX1 NOT_3799 (.Y(I6531),.A(g3186));
INVX1 NOT_3800 (.Y(I11348),.A(g6695));
INVX1 NOT_3801 (.Y(I12344),.A(g7062));
INVX1 NOT_3802 (.Y(I13083),.A(g7921));
INVX1 NOT_3803 (.Y(g3479),.A(g2655));
INVX1 NOT_3804 (.Y(g11195),.A(g11112));
INVX1 NOT_3805 (.Y(g11489),.A(I17482));
INVX1 NOT_3806 (.Y(g6131),.A(g5548));
INVX1 NOT_3807 (.Y(g5661),.A(I9144));
INVX1 NOT_3808 (.Y(g10747),.A(I16432));
INVX1 NOT_3809 (.Y(I15559),.A(g10094));
INVX1 NOT_3810 (.Y(g5075),.A(g4439));
INVX1 NOT_3811 (.Y(g8513),.A(I13708));
INVX1 NOT_3812 (.Y(I15488),.A(g10116));
INVX1 NOT_3813 (.Y(I15424),.A(g10080));
INVX1 NOT_3814 (.Y(g6406),.A(I10314));
INVX1 NOT_3815 (.Y(g10242),.A(I15632));
INVX1 NOT_3816 (.Y(I8007),.A(g3829));
INVX1 NOT_3817 (.Y(g5475),.A(I8892));
INVX1 NOT_3818 (.Y(g4762),.A(I8116));
INVX1 NOT_3819 (.Y(g2798),.A(g2449));
INVX1 NOT_3820 (.Y(g5949),.A(I9591));
INVX1 NOT_3821 (.Y(g7349),.A(I11695));
INVX1 NOT_3822 (.Y(I10192),.A(g6115));
INVX1 NOT_3823 (.Y(g11424),.A(I17327));
INVX1 NOT_3824 (.Y(I9240),.A(g5069));
INVX1 NOT_3825 (.Y(g6635),.A(I10592));
INVX1 NOT_3826 (.Y(I11566),.A(g6820));
INVX1 NOT_3827 (.Y(g11016),.A(I16739));
INVX1 NOT_3828 (.Y(g9108),.A(I14449));
INVX1 NOT_3829 (.Y(g3390),.A(g3161));
INVX1 NOT_3830 (.Y(g9308),.A(I14499));
INVX1 NOT_3831 (.Y(g8036),.A(I12878));
INVX1 NOT_3832 (.Y(g2560),.A(I5684));
INVX1 NOT_3833 (.Y(g5627),.A(g4840));
INVX1 NOT_3834 (.Y(g8436),.A(I13606));
INVX1 NOT_3835 (.Y(g8178),.A(I13083));
INVX1 NOT_3836 (.Y(g6801),.A(I10813));
INVX1 NOT_3837 (.Y(g6305),.A(I10174));
INVX1 NOT_3838 (.Y(I6856),.A(g3318));
INVX1 NOT_3839 (.Y(g4590),.A(I7999));
INVX1 NOT_3840 (.Y(g7848),.A(I12641));
INVX1 NOT_3841 (.Y(g5292),.A(g4445));
INVX1 NOT_3842 (.Y(I10663),.A(g6040));
INVX1 NOT_3843 (.Y(g8378),.A(I13482));
INVX1 NOT_3844 (.Y(g9883),.A(I15060));
INVX1 NOT_3845 (.Y(I9043),.A(g4786));
INVX1 NOT_3846 (.Y(g3501),.A(g3077));
INVX1 NOT_3847 (.Y(I14522),.A(g9108));
INVX1 NOT_3848 (.Y(I8535),.A(g4340));
INVX1 NOT_3849 (.Y(I9443),.A(g5557));
INVX1 NOT_3850 (.Y(g7747),.A(I12406));
INVX1 NOT_3851 (.Y(g5998),.A(I9620));
INVX1 NOT_3852 (.Y(g5646),.A(I9099));
INVX1 NOT_3853 (.Y(g10974),.A(I16723));
INVX1 NOT_3854 (.Y(g8335),.A(I13385));
INVX1 NOT_3855 (.Y(g2873),.A(I6019));
INVX1 NOT_3856 (.Y(g6748),.A(I10753));
INVX1 NOT_3857 (.Y(g2632),.A(g2002));
INVX1 NOT_3858 (.Y(I6074),.A(g2228));
INVX1 NOT_3859 (.Y(g2095),.A(g143));
INVX1 NOT_3860 (.Y(I11653),.A(g6954));
INVX1 NOT_3861 (.Y(g2037),.A(g1771));
INVX1 NOT_3862 (.Y(g8182),.A(I13099));
INVX1 NOT_3863 (.Y(I4886),.A(g257));
INVX1 NOT_3864 (.Y(g4222),.A(g3638));
INVX1 NOT_3865 (.Y(g5603),.A(I9029));
INVX1 NOT_3866 (.Y(I6474),.A(g2297));
INVX1 NOT_3867 (.Y(I7625),.A(g4164));
INVX1 NOT_3868 (.Y(g5039),.A(I8418));
INVX1 NOT_3869 (.Y(I4951),.A(g262));
INVX1 NOT_3870 (.Y(g10293),.A(I15701));
INVX1 NOT_3871 (.Y(g2653),.A(g2011));
INVX1 NOT_3872 (.Y(g2208),.A(g84));
INVX1 NOT_3873 (.Y(g2302),.A(g29));
INVX1 NOT_3874 (.Y(I12029),.A(g6922));
INVX1 NOT_3875 (.Y(g5850),.A(g5320));
INVX1 NOT_3876 (.Y(g6226),.A(I9973));
INVX1 NOT_3877 (.Y(I10553),.A(g6192));
INVX1 NOT_3878 (.Y(g3704),.A(I6861));
INVX1 NOT_3879 (.Y(g8805),.A(I14136));
INVX1 NOT_3880 (.Y(g10265),.A(g10143));
INVX1 NOT_3881 (.Y(g2579),.A(g1969));
INVX1 NOT_3882 (.Y(I5837),.A(g2507));
INVX1 NOT_3883 (.Y(I7938),.A(g3406));
INVX1 NOT_3884 (.Y(I9147),.A(g5011));
INVX1 NOT_3885 (.Y(I13636),.A(g8357));
INVX1 NOT_3886 (.Y(g8422),.A(I13580));
INVX1 NOT_3887 (.Y(I10949),.A(g6747));
INVX1 NOT_3888 (.Y(I17302),.A(g11391));
INVX1 NOT_3889 (.Y(g4899),.A(I8262));
INVX1 NOT_3890 (.Y(I11333),.A(g6670));
INVX1 NOT_3891 (.Y(I13415),.A(g8144));
INVX1 NOT_3892 (.Y(g4464),.A(I7829));
INVX1 NOT_3893 (.Y(g2719),.A(g2043));
INVX1 NOT_3894 (.Y(g9448),.A(g9091));
INVX1 NOT_3895 (.Y(I7909),.A(g3387));
INVX1 NOT_3896 (.Y(I6080),.A(g2108));
INVX1 NOT_3897 (.Y(I14326),.A(g8818));
INVX1 NOT_3898 (.Y(g4785),.A(g3337));
INVX1 NOT_3899 (.Y(g11042),.A(I16787));
INVX1 NOT_3900 (.Y(g10391),.A(g10313));
INVX1 NOT_3901 (.Y(I6480),.A(g2462));
INVX1 NOT_3902 (.Y(g5702),.A(I9243));
INVX1 NOT_3903 (.Y(g6445),.A(I10367));
INVX1 NOT_3904 (.Y(g2752),.A(I5824));
INVX1 NOT_3905 (.Y(I14040),.A(g8649));
INVX1 NOT_3906 (.Y(I14948),.A(g9555));
INVX1 NOT_3907 (.Y(g9827),.A(I14982));
INVX1 NOT_3908 (.Y(g6091),.A(I9744));
INVX1 NOT_3909 (.Y(I10702),.A(g6071));
INVX1 NOT_3910 (.Y(g3810),.A(g3228));
INVX1 NOT_3911 (.Y(g3363),.A(I6549));
INVX1 NOT_3912 (.Y(I10904),.A(g6558));
INVX1 NOT_3913 (.Y(g8798),.A(I14119));
INVX1 NOT_3914 (.Y(g7119),.A(I11354));
INVX1 NOT_3915 (.Y(g7319),.A(I11605));
INVX1 NOT_3916 (.Y(g3432),.A(g3144));
INVX1 NOT_3917 (.Y(I6569),.A(g3186));
INVX1 NOT_3918 (.Y(g10579),.A(g10528));
INVX1 NOT_3919 (.Y(g4563),.A(g3946));
INVX1 NOT_3920 (.Y(g9774),.A(g9474));
INVX1 NOT_3921 (.Y(I7606),.A(g4166));
INVX1 NOT_3922 (.Y(g8560),.A(I13773));
INVX1 NOT_3923 (.Y(I14252),.A(g8783));
INVX1 NOT_3924 (.Y(g6169),.A(I9896));
INVX1 NOT_3925 (.Y(I15383),.A(g10107));
INVX1 NOT_3926 (.Y(I16277),.A(g10536));
INVX1 NOT_3927 (.Y(g6283),.A(I10108));
INVX1 NOT_3928 (.Y(g7352),.A(I11704));
INVX1 NOT_3929 (.Y(g2042),.A(g1796));
INVX1 NOT_3930 (.Y(g4295),.A(I7556));
INVX1 NOT_3931 (.Y(g10578),.A(g10527));
INVX1 NOT_3932 (.Y(I9013),.A(g4767));
INVX1 NOT_3933 (.Y(g4237),.A(g4013));
INVX1 NOT_3934 (.Y(g6407),.A(I10317));
INVX1 NOT_3935 (.Y(I14564),.A(g9026));
INVX1 NOT_3936 (.Y(g6920),.A(I11034));
INVX1 NOT_3937 (.Y(g6578),.A(I10526));
INVX1 NOT_3938 (.Y(g6868),.A(I10946));
INVX1 NOT_3939 (.Y(g5616),.A(I9046));
INVX1 NOT_3940 (.Y(I16595),.A(g10783));
INVX1 NOT_3941 (.Y(g8873),.A(I14191));
INVX1 NOT_3942 (.Y(g8632),.A(I13915));
INVX1 NOT_3943 (.Y(g8095),.A(g7942));
INVX1 NOT_3944 (.Y(g2164),.A(I5095));
INVX1 NOT_3945 (.Y(g6718),.A(g5949));
INVX1 NOT_3946 (.Y(g2364),.A(g611));
INVX1 NOT_3947 (.Y(g2233),.A(I5224));
INVX1 NOT_3948 (.Y(g9780),.A(g9474));
INVX1 NOT_3949 (.Y(g4194),.A(I7399));
INVX1 NOT_3950 (.Y(I16623),.A(g10858));
INVX1 NOT_3951 (.Y(g8437),.A(I13609));
INVX1 NOT_3952 (.Y(I10183),.A(g6108));
INVX1 NOT_3953 (.Y(I7586),.A(g4127));
INVX1 NOT_3954 (.Y(g11065),.A(g10974));
INVX1 NOT_3955 (.Y(g4394),.A(I7729));
INVX1 NOT_3956 (.Y(I5192),.A(g55));
INVX1 NOT_3957 (.Y(I6976),.A(g2884));
INVX1 NOT_3958 (.Y(g2054),.A(g1864));
INVX1 NOT_3959 (.Y(g6582),.A(g5949));
INVX1 NOT_3960 (.Y(I13609),.A(g8312));
INVX1 NOT_3961 (.Y(I14397),.A(g8888));
INVX1 NOT_3962 (.Y(g7386),.A(I11767));
INVX1 NOT_3963 (.Y(g4731),.A(I8085));
INVX1 NOT_3964 (.Y(I11312),.A(g6488));
INVX1 NOT_3965 (.Y(g5647),.A(I9102));
INVX1 NOT_3966 (.Y(g2454),.A(I5549));
INVX1 NOT_3967 (.Y(g8579),.A(I13822));
INVX1 NOT_3968 (.Y(g8869),.A(I14179));
INVX1 NOT_3969 (.Y(g7975),.A(I12773));
INVX1 NOT_3970 (.Y(I13200),.A(g8251));
INVX1 NOT_3971 (.Y(g6261),.A(I10042));
INVX1 NOT_3972 (.Y(I11608),.A(g6903));
INVX1 NOT_3973 (.Y(g2296),.A(I5332));
INVX1 NOT_3974 (.Y(I11115),.A(g6462));
INVX1 NOT_3975 (.Y(I12604),.A(g7630));
INVX1 NOT_3976 (.Y(g10116),.A(I15356));
INVX1 NOT_3977 (.Y(I9117),.A(g5615));
INVX1 NOT_3978 (.Y(g6793),.A(I10795));
INVX1 NOT_3979 (.Y(g8719),.A(g8579));
INVX1 NOT_3980 (.Y(g4557),.A(g3946));
INVX1 NOT_3981 (.Y(I9317),.A(g5576));
INVX1 NOT_3982 (.Y(g2725),.A(g2018));
INVX1 NOT_3983 (.Y(g1974),.A(g627));
INVX1 NOT_3984 (.Y(I14509),.A(g8926));
INVX1 NOT_3985 (.Y(g5546),.A(I8973));
INVX1 NOT_3986 (.Y(g7026),.A(I11173));
INVX1 NOT_3987 (.Y(I5854),.A(g2523));
INVX1 NOT_3988 (.Y(I8388),.A(g4239));
INVX1 NOT_3989 (.Y(g4966),.A(I8340));
INVX1 NOT_3990 (.Y(I12770),.A(g7638));
INVX1 NOT_3991 (.Y(I14933),.A(g9454));
INVX1 NOT_3992 (.Y(g7426),.A(I11814));
INVX1 NOT_3993 (.Y(g9994),.A(I15196));
INVX1 NOT_3994 (.Y(g9290),.A(I14494));
INVX1 NOT_3995 (.Y(I11921),.A(g6904));
INVX1 NOT_3996 (.Y(I17662),.A(g11602));
INVX1 NOT_3997 (.Y(I12981),.A(g8041));
INVX1 NOT_3998 (.Y(g8752),.A(g8635));
INVX1 NOT_3999 (.Y(g6227),.A(g5446));
INVX1 NOT_4000 (.Y(g10041),.A(I15250));
INVX1 NOT_4001 (.Y(g5503),.A(g4515));
INVX1 NOT_4002 (.Y(I7710),.A(g3749));
INVX1 NOT_4003 (.Y(g7614),.A(I12190));
INVX1 NOT_4004 (.Y(g10275),.A(I15669));
INVX1 NOT_4005 (.Y(g4242),.A(g3664));
INVX1 NOT_4006 (.Y(g10493),.A(I16114));
INVX1 NOT_4007 (.Y(g7325),.A(I11623));
INVX1 NOT_4008 (.Y(I17249),.A(g11342));
INVX1 NOT_4009 (.Y(g4948),.A(I8315));
INVX1 NOT_4010 (.Y(I7691),.A(g3363));
INVX1 NOT_4011 (.Y(g9816),.A(g9490));
INVX1 NOT_4012 (.Y(I17482),.A(g11479));
INVX1 NOT_4013 (.Y(g10465),.A(I15986));
INVX1 NOT_4014 (.Y(g1980),.A(g646));
INVX1 NOT_4015 (.Y(I8247),.A(g4615));
INVX1 NOT_4016 (.Y(g7984),.A(I12796));
INVX1 NOT_4017 (.Y(g2012),.A(g981));
INVX1 NOT_4018 (.Y(g11160),.A(g10950));
INVX1 NOT_4019 (.Y(g8442),.A(I13624));
INVX1 NOT_4020 (.Y(I17710),.A(g11620));
INVX1 NOT_4021 (.Y(g6203),.A(g5446));
INVX1 NOT_4022 (.Y(I17552),.A(g11502));
INVX1 NOT_4023 (.Y(I16853),.A(g10907));
INVX1 NOT_4024 (.Y(I9581),.A(g5111));
INVX1 NOT_4025 (.Y(g10035),.A(I15241));
INVX1 NOT_4026 (.Y(g5120),.A(I8520));
INVX1 NOT_4027 (.Y(I5031),.A(g928));
INVX1 NOT_4028 (.Y(g5320),.A(g4418));
INVX1 NOT_4029 (.Y(g4254),.A(g4013));
INVX1 NOT_4030 (.Y(I16589),.A(g10820));
INVX1 NOT_4031 (.Y(I11674),.A(g7051));
INVX1 NOT_4032 (.Y(g10806),.A(I16518));
INVX1 NOT_4033 (.Y(g7544),.A(I11964));
INVX1 NOT_4034 (.Y(g8164),.A(g7872));
INVX1 NOT_4035 (.Y(I13674),.A(g8304));
INVX1 NOT_4036 (.Y(I15470),.A(g10111));
INVX1 NOT_4037 (.Y(I5812),.A(g2090));
INVX1 NOT_4038 (.Y(g8233),.A(g7872));
INVX1 NOT_4039 (.Y(g11617),.A(I17669));
INVX1 NOT_4040 (.Y(I6183),.A(g2131));
INVX1 NOT_4041 (.Y(g11470),.A(I17447));
INVX1 NOT_4042 (.Y(I7659),.A(g3731));
INVX1 NOT_4043 (.Y(g10142),.A(I15424));
INVX1 NOT_4044 (.Y(g2888),.A(I6046));
INVX1 NOT_4045 (.Y(I6924),.A(g2843));
INVX1 NOT_4046 (.Y(g7636),.A(I12248));
INVX1 NOT_4047 (.Y(I6220),.A(g883));
INVX1 NOT_4048 (.Y(I4891),.A(g582));
INVX1 NOT_4049 (.Y(g2171),.A(I5116));
INVX1 NOT_4050 (.Y(g4438),.A(I7790));
INVX1 NOT_4051 (.Y(I14452),.A(g8922));
INVX1 NOT_4052 (.Y(g4773),.A(I8133));
INVX1 NOT_4053 (.Y(g7306),.A(I11566));
INVX1 NOT_4054 (.Y(I13732),.A(g8291));
INVX1 NOT_4055 (.Y(g8296),.A(I13242));
INVX1 NOT_4056 (.Y(g2956),.A(I6159));
INVX1 NOT_4057 (.Y(I15075),.A(g9761));
INVX1 NOT_4058 (.Y(g8725),.A(g8589));
INVX1 NOT_4059 (.Y(g7790),.A(I12535));
INVX1 NOT_4060 (.Y(g9263),.A(g8892));
INVX1 NOT_4061 (.Y(g3683),.A(I6844));
INVX1 NOT_4062 (.Y(g11075),.A(g10937));
INVX1 NOT_4063 (.Y(I5765),.A(g2004));
INVX1 NOT_4064 (.Y(I15595),.A(g10165));
INVX1 NOT_4065 (.Y(I15467),.A(g10079));
INVX1 NOT_4066 (.Y(I15494),.A(g10117));
INVX1 NOT_4067 (.Y(I17356),.A(g11384));
INVX1 NOT_4068 (.Y(g8532),.A(I13741));
INVX1 NOT_4069 (.Y(I8308),.A(g4443));
INVX1 NOT_4070 (.Y(g7187),.A(I11405));
INVX1 NOT_4071 (.Y(I7311),.A(g2803));
INVX1 NOT_4072 (.Y(g4769),.A(g3586));
INVX1 NOT_4073 (.Y(g5987),.A(I9605));
INVX1 NOT_4074 (.Y(I11692),.A(g7048));
INVX1 NOT_4075 (.Y(g7387),.A(I11770));
INVX1 NOT_4076 (.Y(g11467),.A(I17438));
INVX1 NOT_4077 (.Y(I9995),.A(g5536));
INVX1 NOT_4078 (.Y(I12832),.A(g7681));
INVX1 NOT_4079 (.Y(I4859),.A(g578));
INVX1 NOT_4080 (.Y(I10051),.A(g5702));
INVX1 NOT_4081 (.Y(I10072),.A(g5719));
INVX1 NOT_4082 (.Y(g4212),.A(I7453));
INVX1 NOT_4083 (.Y(I9479),.A(g4954));
INVX1 NOT_4084 (.Y(g6689),.A(g5830));
INVX1 NOT_4085 (.Y(g10130),.A(I15392));
INVX1 NOT_4086 (.Y(g7756),.A(I12433));
INVX1 NOT_4087 (.Y(g2297),.A(g865));
INVX1 NOT_4088 (.Y(g11623),.A(I17687));
INVX1 NOT_4089 (.Y(g6388),.A(I10286));
INVX1 NOT_4090 (.Y(g10193),.A(g10057));
INVX1 NOT_4091 (.Y(I16616),.A(g10796));
INVX1 NOT_4092 (.Y(g11037),.A(I16772));
INVX1 NOT_4093 (.Y(I10592),.A(g5865));
INVX1 NOT_4094 (.Y(g5299),.A(g4393));
INVX1 NOT_4095 (.Y(I10756),.A(g5810));
INVX1 NOT_4096 (.Y(I15782),.A(g10259));
INVX1 NOT_4097 (.Y(g7622),.A(g7067));
INVX1 NOT_4098 (.Y(g3735),.A(I6921));
INVX1 NOT_4099 (.Y(g7027),.A(I11176));
INVX1 NOT_4100 (.Y(g7427),.A(I11817));
INVX1 NOT_4101 (.Y(I17182),.A(g11309));
INVX1 NOT_4102 (.Y(g10165),.A(I15491));
INVX1 NOT_4103 (.Y(I13400),.A(g8236));
INVX1 NOT_4104 (.Y(g10523),.A(g10456));
INVX1 NOT_4105 (.Y(I17672),.A(g11605));
INVX1 NOT_4106 (.Y(g3782),.A(I7006));
INVX1 NOT_4107 (.Y(I13013),.A(g8048));
INVX1 NOT_4108 (.Y(g5892),.A(I9519));
INVX1 NOT_4109 (.Y(I11214),.A(g6528));
INVX1 NOT_4110 (.Y(g7904),.A(I12690));
INVX1 NOT_4111 (.Y(g11419),.A(I17312));
INVX1 NOT_4112 (.Y(g2745),.A(I5809));
INVX1 NOT_4113 (.Y(g2639),.A(I5754));
INVX1 NOT_4114 (.Y(g6030),.A(I9639));
INVX1 NOT_4115 (.Y(g2338),.A(g1909));
INVX1 NOT_4116 (.Y(g11352),.A(I17173));
INVX1 NOT_4117 (.Y(I15418),.A(g10083));
INVX1 NOT_4118 (.Y(I5073),.A(g34));
INVX1 NOT_4119 (.Y(I13329),.A(g8116));
INVX1 NOT_4120 (.Y(I11207),.A(g6524));
INVX1 NOT_4121 (.Y(g7446),.A(g7148));
INVX1 NOT_4122 (.Y(g3475),.A(g3056));
INVX1 NOT_4123 (.Y(I6999),.A(g2905));
INVX1 NOT_4124 (.Y(g11155),.A(g10950));
INVX1 NOT_4125 (.Y(I7284),.A(g3255));
INVX1 NOT_4126 (.Y(I15266),.A(g10001));
INVX1 NOT_4127 (.Y(g8990),.A(I14391));
INVX1 NOT_4128 (.Y(I9156),.A(g5032));
INVX1 NOT_4129 (.Y(I12099),.A(g7258));
INVX1 NOT_4130 (.Y(I11005),.A(g6386));
INVX1 NOT_4131 (.Y(I12388),.A(g7219));
INVX1 NOT_4132 (.Y(I17331),.A(g11357));
INVX1 NOT_4133 (.Y(I13005),.A(g8046));
INVX1 NOT_4134 (.Y(g8888),.A(I14232));
INVX1 NOT_4135 (.Y(g7403),.A(I11783));
INVX1 NOT_4136 (.Y(g3627),.A(I6784));
INVX1 NOT_4137 (.Y(g4822),.A(g3706));
INVX1 NOT_4138 (.Y(g8029),.A(I12871));
INVX1 NOT_4139 (.Y(g6564),.A(g5784));
INVX1 NOT_4140 (.Y(I16808),.A(g10906));
INVX1 NOT_4141 (.Y(g8171),.A(I13068));
INVX1 NOT_4142 (.Y(g7345),.A(I11683));
INVX1 NOT_4143 (.Y(I17513),.A(g11482));
INVX1 NOT_4144 (.Y(I8711),.A(g4530));
INVX1 NOT_4145 (.Y(g2808),.A(g2156));
INVX1 NOT_4146 (.Y(g3292),.A(g2373));
INVX1 NOT_4147 (.Y(I10846),.A(g6729));
INVX1 NOT_4148 (.Y(g8787),.A(I14094));
INVX1 NOT_4149 (.Y(I12251),.A(g7076));
INVX1 NOT_4150 (.Y(g7763),.A(I12454));
INVX1 NOT_4151 (.Y(I16101),.A(g10381));
INVX1 NOT_4152 (.Y(g8956),.A(I14319));
INVX1 NOT_4153 (.Y(g2707),.A(g2041));
INVX1 NOT_4154 (.Y(I8827),.A(g4477));
INVX1 NOT_4155 (.Y(g10437),.A(g10333));
INVX1 NOT_4156 (.Y(I8133),.A(g3632));
INVX1 NOT_4157 (.Y(g2759),.A(I5843));
INVX1 NOT_4158 (.Y(I8333),.A(g4456));
INVX1 NOT_4159 (.Y(I7420),.A(g4167));
INVX1 NOT_4160 (.Y(g7637),.A(I12251));
INVX1 NOT_4161 (.Y(I15589),.A(g10161));
INVX1 NOT_4162 (.Y(g5078),.A(g4372));
INVX1 NOT_4163 (.Y(g3039),.A(g2310));
INVX1 NOT_4164 (.Y(g2201),.A(g102));
INVX1 NOT_4165 (.Y(g3439),.A(g3144));
INVX1 NOT_4166 (.Y(g7107),.A(I11342));
INVX1 NOT_4167 (.Y(I7559),.A(g4116));
INVX1 NOT_4168 (.Y(g7307),.A(I11569));
INVX1 NOT_4169 (.Y(I12032),.A(g6923));
INVX1 NOT_4170 (.Y(g8297),.A(I13245));
INVX1 NOT_4171 (.Y(g10347),.A(I15807));
INVX1 NOT_4172 (.Y(g5035),.A(I8410));
INVX1 NOT_4173 (.Y(I6944),.A(g2859));
INVX1 NOT_4174 (.Y(I8396),.A(g4255));
INVX1 NOT_4175 (.Y(g10253),.A(g10138));
INVX1 NOT_4176 (.Y(I6240),.A(g878));
INVX1 NOT_4177 (.Y(I7931),.A(g3624));
INVX1 NOT_4178 (.Y(g7359),.A(I11725));
INVX1 NOT_4179 (.Y(g6108),.A(I9779));
INVX1 NOT_4180 (.Y(g6308),.A(I10183));
INVX1 NOT_4181 (.Y(I9810),.A(g5576));
INVX1 NOT_4182 (.Y(g5082),.A(g4840));
INVX1 NOT_4183 (.Y(g2449),.A(g790));
INVX1 NOT_4184 (.Y(I9032),.A(g4732));
INVX1 NOT_4185 (.Y(I11100),.A(g6442));
INVX1 NOT_4186 (.Y(g5482),.A(I8903));
INVX1 NOT_4187 (.Y(I14405),.A(g8937));
INVX1 NOT_4188 (.Y(g10600),.A(I16277));
INVX1 NOT_4189 (.Y(g11401),.A(I17246));
INVX1 NOT_4190 (.Y(g10781),.A(I16475));
INVX1 NOT_4191 (.Y(I4783),.A(g873));
INVX1 NOT_4192 (.Y(I6043),.A(g2267));
INVX1 NOT_4193 (.Y(I9053),.A(g4752));
INVX1 NOT_4194 (.Y(g8684),.A(I13969));
INVX1 NOT_4195 (.Y(g3583),.A(I6742));
INVX1 NOT_4196 (.Y(g4895),.A(I8250));
INVX1 NOT_4197 (.Y(g5876),.A(g5361));
INVX1 NOT_4198 (.Y(g8138),.A(I13013));
INVX1 NOT_4199 (.Y(I6443),.A(g2363));
INVX1 NOT_4200 (.Y(I11235),.A(g6538));
INVX1 NOT_4201 (.Y(g8338),.A(I13394));
INVX1 NOT_4202 (.Y(g10236),.A(g10190));
INVX1 NOT_4203 (.Y(g7757),.A(I12436));
INVX1 NOT_4204 (.Y(g2604),.A(I5713));
INVX1 NOT_4205 (.Y(g4062),.A(I7185));
INVX1 NOT_4206 (.Y(g2098),.A(I4938));
INVX1 NOT_4207 (.Y(I11683),.A(g7069));
INVX1 NOT_4208 (.Y(g5656),.A(I9129));
INVX1 NOT_4209 (.Y(g7416),.A(I11800));
INVX1 NOT_4210 (.Y(g4620),.A(I8031));
INVX1 NOT_4211 (.Y(g10351),.A(I15817));
INVX1 NOT_4212 (.Y(g4462),.A(I7825));
INVX1 NOT_4213 (.Y(I15864),.A(g10339));
INVX1 NOT_4214 (.Y(I5399),.A(g895));
INVX1 NOT_4215 (.Y(g6589),.A(I10549));
INVX1 NOT_4216 (.Y(I12871),.A(g7638));
INVX1 NOT_4217 (.Y(g10175),.A(I15517));
INVX1 NOT_4218 (.Y(g10821),.A(I16531));
INVX1 NOT_4219 (.Y(I7630),.A(g3524));
INVX1 NOT_4220 (.Y(I15749),.A(g10263));
INVX1 NOT_4221 (.Y(g2833),.A(I5949));
INVX1 NOT_4222 (.Y(I6034),.A(g2210));
INVX1 NOT_4223 (.Y(g7522),.A(I11904));
INVX1 NOT_4224 (.Y(I8418),.A(g4794));
INVX1 NOT_4225 (.Y(g7811),.A(I12598));
INVX1 NOT_4226 (.Y(g7315),.A(I11593));
INVX1 NOT_4227 (.Y(g11616),.A(I17666));
INVX1 NOT_4228 (.Y(I17149),.A(g11306));
INVX1 NOT_4229 (.Y(I6565),.A(g2614));
INVX1 NOT_4230 (.Y(g7047),.A(I11222));
INVX1 NOT_4231 (.Y(I7300),.A(g2883));
INVX1 NOT_4232 (.Y(g11313),.A(I17104));
INVX1 NOT_4233 (.Y(I12360),.A(g7183));
INVX1 NOT_4234 (.Y(I8290),.A(g4778));
INVX1 NOT_4235 (.Y(g10063),.A(I15287));
INVX1 NOT_4236 (.Y(I17387),.A(g11438));
INVX1 NOT_4237 (.Y(g8707),.A(g8671));
INVX1 NOT_4238 (.Y(g6165),.A(g5446));
INVX1 NOT_4239 (.Y(g10264),.A(g10128));
INVX1 NOT_4240 (.Y(g6571),.A(I10503));
INVX1 NOT_4241 (.Y(g6365),.A(I10274));
INVX1 NOT_4242 (.Y(g6861),.A(I10941));
INVX1 NOT_4243 (.Y(g5214),.A(g4640));
INVX1 NOT_4244 (.Y(g10137),.A(I15409));
INVX1 NOT_4245 (.Y(g6048),.A(I9673));
INVX1 NOT_4246 (.Y(I11515),.A(g6589));
INVX1 NOT_4247 (.Y(g9772),.A(g9432));
INVX1 NOT_4248 (.Y(I11882),.A(g6895));
INVX1 NOT_4249 (.Y(I5510),.A(g588));
INVX1 NOT_4250 (.Y(g2539),.A(I5652));
INVX1 NOT_4251 (.Y(g2896),.A(g2356));
INVX1 NOT_4252 (.Y(I6347),.A(g2462));
INVX1 NOT_4253 (.Y(I15704),.A(g10238));
INVX1 NOT_4254 (.Y(I5245),.A(g925));
INVX1 NOT_4255 (.Y(g6448),.A(I10374));
INVX1 NOT_4256 (.Y(g9531),.A(I14678));
INVX1 NOT_4257 (.Y(I15305),.A(g10001));
INVX1 NOT_4258 (.Y(g6711),.A(g5949));
INVX1 NOT_4259 (.Y(g6055),.A(I9688));
INVX1 NOT_4260 (.Y(I12162),.A(g7146));
INVX1 NOT_4261 (.Y(I17104),.A(g11223));
INVX1 NOT_4262 (.Y(g10873),.A(I16589));
INVX1 NOT_4263 (.Y(g11053),.A(g10950));
INVX1 NOT_4264 (.Y(I8256),.A(g4711));
INVX1 NOT_4265 (.Y(g9890),.A(I15075));
INVX1 NOT_4266 (.Y(I10282),.A(g6163));
INVX1 NOT_4267 (.Y(g3404),.A(g3121));
INVX1 NOT_4268 (.Y(g6133),.A(I9836));
INVX1 NOT_4269 (.Y(g11466),.A(I17435));
INVX1 NOT_4270 (.Y(g5663),.A(I9150));
INVX1 NOT_4271 (.Y(I10302),.A(g6179));
INVX1 NOT_4272 (.Y(I6914),.A(g2828));
INVX1 NOT_4273 (.Y(g9505),.A(g9052));
INVX1 NOT_4274 (.Y(g2162),.A(I5089));
INVX1 NOT_4275 (.Y(I7973),.A(g3437));
INVX1 NOT_4276 (.Y(I15036),.A(g9721));
INVX1 NOT_4277 (.Y(g2268),.A(g654));
INVX1 NOT_4278 (.Y(g8449),.A(I13645));
INVX1 NOT_4279 (.Y(g4192),.A(I7393));
INVX1 NOT_4280 (.Y(I10105),.A(g5736));
INVX1 NOT_4281 (.Y(g4298),.A(g4130));
INVX1 NOT_4282 (.Y(g3764),.A(I6971));
INVX1 NOT_4283 (.Y(I12451),.A(g7538));
INVX1 NOT_4284 (.Y(g6846),.A(I10910));
INVX1 NOT_4285 (.Y(g11036),.A(I16769));
INVX1 NOT_4286 (.Y(I12472),.A(g7539));
INVX1 NOT_4287 (.Y(g8575),.A(I13816));
INVX1 NOT_4288 (.Y(g3546),.A(g3307));
INVX1 NOT_4289 (.Y(I14105),.A(g8776));
INVX1 NOT_4290 (.Y(g4485),.A(g3546));
INVX1 NOT_4291 (.Y(I6013),.A(g2200));
INVX1 NOT_4292 (.Y(g5402),.A(I8842));
INVX1 NOT_4293 (.Y(g6196),.A(g5446));
INVX1 NOT_4294 (.Y(g7880),.A(g7479));
INVX1 NOT_4295 (.Y(g6396),.A(I10296));
INVX1 NOT_4296 (.Y(g7595),.A(I12123));
INVX1 NOT_4297 (.Y(g6803),.A(I10819));
INVX1 NOT_4298 (.Y(g7537),.A(I11947));
INVX1 NOT_4299 (.Y(g5236),.A(g4361));
INVX1 NOT_4300 (.Y(I17368),.A(g11423));
INVX1 NOT_4301 (.Y(g8604),.A(g8479));
INVX1 NOT_4302 (.Y(g10208),.A(I15580));
INVX1 NOT_4303 (.Y(I16239),.A(g10525));
INVX1 NOT_4304 (.Y(g11642),.A(I17730));
INVX1 NOT_4305 (.Y(g8498),.A(g8353));
INVX1 NOT_4306 (.Y(I11584),.A(g6827));
INVX1 NOT_4307 (.Y(g1972),.A(g461));
INVX1 NOT_4308 (.Y(I8421),.A(g4309));
INVX1 NOT_4309 (.Y(g9474),.A(g9331));
INVX1 NOT_4310 (.Y(g7272),.A(I11519));
INVX1 NOT_4311 (.Y(I13206),.A(g8197));
INVX1 NOT_4312 (.Y(g10542),.A(I16193));
INVX1 NOT_4313 (.Y(g6509),.A(I10427));
INVX1 NOT_4314 (.Y(g11064),.A(g10974));
INVX1 NOT_4315 (.Y(I15733),.A(g10257));
INVX1 NOT_4316 (.Y(g7612),.A(I12186));
INVX1 NOT_4317 (.Y(g7243),.A(I11483));
INVX1 NOT_4318 (.Y(g2086),.A(I4906));
INVX1 NOT_4319 (.Y(I11759),.A(g7244));
INVX1 NOT_4320 (.Y(I11725),.A(g7040));
INVX1 NOT_4321 (.Y(I12776),.A(g7586));
INVX1 NOT_4322 (.Y(g5657),.A(I9132));
INVX1 NOT_4323 (.Y(g10913),.A(I16691));
INVX1 NOT_4324 (.Y(I16941),.A(g11076));
INVX1 NOT_4325 (.Y(g2728),.A(g2025));
INVX1 NOT_4326 (.Y(I13114),.A(g7930));
INVX1 NOT_4327 (.Y(g6418),.A(g6137));
INVX1 NOT_4328 (.Y(I11082),.A(g6749));
INVX1 NOT_4329 (.Y(g7982),.A(I12790));
INVX1 NOT_4330 (.Y(g4520),.A(I7923));
INVX1 NOT_4331 (.Y(g5222),.A(g4640));
INVX1 NOT_4332 (.Y(I17228),.A(g11300));
INVX1 NOT_4333 (.Y(g11630),.A(I17704));
INVX1 NOT_4334 (.Y(g2185),.A(g46));
INVX1 NOT_4335 (.Y(g4219),.A(g3635));
INVX1 NOT_4336 (.Y(g6290),.A(I10129));
INVX1 NOT_4337 (.Y(I7151),.A(g2642));
INVX1 NOT_4338 (.Y(g2881),.A(I6031));
INVX1 NOT_4339 (.Y(I7351),.A(g4061));
INVX1 NOT_4340 (.Y(I16518),.A(g10718));
INVX1 NOT_4341 (.Y(I6601),.A(g3186));
INVX1 NOT_4342 (.Y(I7648),.A(g3727));
INVX1 NOT_4343 (.Y(I12825),.A(g7696));
INVX1 NOT_4344 (.Y(g10320),.A(I15756));
INVX1 NOT_4345 (.Y(g10905),.A(I16667));
INVX1 NOT_4346 (.Y(g7629),.A(I12229));
INVX1 NOT_4347 (.Y(I15665),.A(g10193));
INVX1 NOT_4348 (.Y(g7328),.A(I11632));
INVX1 NOT_4349 (.Y(g2070),.A(g213));
INVX1 NOT_4350 (.Y(g10530),.A(g10466));
INVX1 NOT_4351 (.Y(g3906),.A(g3015));
INVX1 NOT_4352 (.Y(I17716),.A(g11622));
INVX1 NOT_4353 (.Y(g7330),.A(I11638));
INVX1 NOT_4354 (.Y(g10593),.A(I16264));
INVX1 NOT_4355 (.Y(I4866),.A(g579));
INVX1 NOT_4356 (.Y(g8362),.A(I13466));
INVX1 NOT_4357 (.Y(I13744),.A(g8297));
INVX1 NOT_4358 (.Y(g2025),.A(g1696));
INVX1 NOT_4359 (.Y(I11345),.A(g6692));
INVX1 NOT_4360 (.Y(g10346),.A(I15804));
INVX1 NOT_4361 (.Y(I8631),.A(g4425));
INVX1 NOT_4362 (.Y(g5899),.A(g5361));
INVX1 NOT_4363 (.Y(g8419),.A(I13571));
INVX1 NOT_4364 (.Y(g4958),.A(I8328));
INVX1 NOT_4365 (.Y(g6256),.A(I10027));
INVX1 NOT_4366 (.Y(g4176),.A(I7345));
INVX1 NOT_4367 (.Y(g6816),.A(I10858));
INVX1 NOT_4368 (.Y(g10122),.A(I15374));
INVX1 NOT_4369 (.Y(g4376),.A(I7691));
INVX1 NOT_4370 (.Y(g4005),.A(I7143));
INVX1 NOT_4371 (.Y(g10464),.A(I15983));
INVX1 NOT_4372 (.Y(I10027),.A(g5751));
INVX1 NOT_4373 (.Y(I15476),.A(g10114));
INVX1 NOT_4374 (.Y(I15485),.A(g10092));
INVX1 NOT_4375 (.Y(g7800),.A(I12565));
INVX1 NOT_4376 (.Y(g10034),.A(I15238));
INVX1 NOT_4377 (.Y(g6181),.A(g5426));
INVX1 NOT_4378 (.Y(I11804),.A(g7190));
INVX1 NOT_4379 (.Y(I14249),.A(g8804));
INVX1 NOT_4380 (.Y(g11454),.A(I17419));
INVX1 NOT_4381 (.Y(g6847),.A(g6482));
INVX1 NOT_4382 (.Y(g10292),.A(I15698));
INVX1 NOT_4383 (.Y(I9475),.A(g5445));
INVX1 NOT_4384 (.Y(I10248),.A(g6125));
INVX1 NOT_4385 (.Y(g6685),.A(I10648));
INVX1 NOT_4386 (.Y(g6197),.A(I9930));
INVX1 NOT_4387 (.Y(g6700),.A(g5949));
INVX1 NOT_4388 (.Y(I17112),.A(g11227));
INVX1 NOT_4389 (.Y(I10710),.A(g6088));
INVX1 NOT_4390 (.Y(g6397),.A(I10299));
INVX1 NOT_4391 (.Y(I10003),.A(g4908));
INVX1 NOT_4392 (.Y(g7213),.A(I11447));
INVX1 NOT_4393 (.Y(I10204),.A(g6031));
INVX1 NOT_4394 (.Y(I14552),.A(g9264));
INVX1 NOT_4395 (.Y(I5336),.A(g1700));
INVX1 NOT_4396 (.Y(g2131),.A(I5060));
INVX1 NOT_4397 (.Y(g8486),.A(g8348));
INVX1 NOT_4398 (.Y(I6784),.A(g2742));
INVX1 NOT_4399 (.Y(g2006),.A(g932));
INVX1 NOT_4400 (.Y(g2331),.A(g658));
INVX1 NOT_4401 (.Y(I16577),.A(g10825));
INVX1 NOT_4402 (.Y(g4733),.A(I8089));
INVX1 NOT_4403 (.Y(g2406),.A(g1365));
INVX1 NOT_4404 (.Y(g5844),.A(I9461));
INVX1 NOT_4405 (.Y(I13332),.A(g8206));
INVX1 NOT_4406 (.Y(g6263),.A(I10048));
INVX1 NOT_4407 (.Y(g4270),.A(g4013));
INVX1 NOT_4408 (.Y(I11135),.A(g6679));
INVX1 NOT_4409 (.Y(I7372),.A(g4057));
INVX1 NOT_4410 (.Y(g10136),.A(I15406));
INVX1 NOT_4411 (.Y(g2635),.A(g2003));
INVX1 NOT_4412 (.Y(I16439),.A(g10702));
INVX1 NOT_4413 (.Y(I17742),.A(g11636));
INVX1 NOT_4414 (.Y(I12318),.A(g6862));
INVX1 NOT_4415 (.Y(g11074),.A(g10901));
INVX1 NOT_4416 (.Y(g6950),.A(I11094));
INVX1 NOT_4417 (.Y(g11239),.A(g11112));
INVX1 NOT_4418 (.Y(I10081),.A(g5735));
INVX1 NOT_4419 (.Y(I17096),.A(g11219));
INVX1 NOT_4420 (.Y(g4225),.A(I7478));
INVX1 NOT_4421 (.Y(I15238),.A(g9974));
INVX1 NOT_4422 (.Y(g2087),.A(g225));
INVX1 NOT_4423 (.Y(g11594),.A(I17636));
INVX1 NOT_4424 (.Y(g3945),.A(I7096));
INVX1 NOT_4425 (.Y(I7143),.A(g2614));
INVX1 NOT_4426 (.Y(I5943),.A(g2233));
INVX1 NOT_4427 (.Y(g2801),.A(g2117));
INVX1 NOT_4428 (.Y(g5089),.A(g4840));
INVX1 NOT_4429 (.Y(I13406),.A(g8179));
INVX1 NOT_4430 (.Y(I9084),.A(g4886));
INVX1 NOT_4431 (.Y(g3738),.A(g3062));
INVX1 NOT_4432 (.Y(I13962),.A(g8451));
INVX1 NOT_4433 (.Y(I14786),.A(g9266));
INVX1 NOT_4434 (.Y(g7512),.A(g7148));
INVX1 NOT_4435 (.Y(g8025),.A(I12867));
INVX1 NOT_4436 (.Y(g9760),.A(g9454));
INVX1 NOT_4437 (.Y(I6294),.A(g2238));
INVX1 NOT_4438 (.Y(I17681),.A(g11608));
INVX1 NOT_4439 (.Y(g8425),.A(I13589));
INVX1 NOT_4440 (.Y(g3709),.A(I6870));
INVX1 NOT_4441 (.Y(g4124),.A(I7269));
INVX1 NOT_4442 (.Y(g4324),.A(g4144));
INVX1 NOT_4443 (.Y(g2748),.A(I5812));
INVX1 NOT_4444 (.Y(g6562),.A(g5774));
INVX1 NOT_4445 (.Y(g7366),.A(I11746));
INVX1 NOT_4446 (.Y(g10164),.A(I15488));
INVX1 NOT_4447 (.Y(I11833),.A(g7077));
INVX1 NOT_4448 (.Y(I11049),.A(g6635));
INVX1 NOT_4449 (.Y(I15675),.A(g10133));
INVX1 NOT_4450 (.Y(g4469),.A(I7840));
INVX1 NOT_4451 (.Y(g5705),.A(I9248));
INVX1 NOT_4452 (.Y(g5471),.A(g4370));
INVX1 NOT_4453 (.Y(g2755),.A(I5833));
INVX1 NOT_4454 (.Y(g11185),.A(I16956));
INVX1 NOT_4455 (.Y(g7056),.A(I11249));
INVX1 NOT_4456 (.Y(I17730),.A(g11638));
INVX1 NOT_4457 (.Y(g3907),.A(I7076));
INVX1 NOT_4458 (.Y(g10891),.A(I16635));
INVX1 NOT_4459 (.Y(g2226),.A(g86));
INVX1 NOT_4460 (.Y(I6501),.A(g2578));
INVX1 NOT_4461 (.Y(I10090),.A(g5767));
INVX1 NOT_4462 (.Y(g6723),.A(I10716));
INVX1 NOT_4463 (.Y(I13048),.A(g8059));
INVX1 NOT_4464 (.Y(g6257),.A(I10030));
INVX1 NOT_4465 (.Y(I14090),.A(g8771));
INVX1 NOT_4466 (.Y(g11518),.A(I17563));
INVX1 NOT_4467 (.Y(g4177),.A(I7348));
INVX1 NOT_4468 (.Y(I6156),.A(g2119));
INVX1 NOT_4469 (.Y(g6101),.A(I9762));
INVX1 NOT_4470 (.Y(g7148),.A(I11397));
INVX1 NOT_4471 (.Y(g6817),.A(I10861));
INVX1 NOT_4472 (.Y(g7649),.A(I12258));
INVX1 NOT_4473 (.Y(g5948),.A(I9588));
INVX1 NOT_4474 (.Y(g6301),.A(I10162));
INVX1 NOT_4475 (.Y(g7348),.A(I11692));
INVX1 NOT_4476 (.Y(I6356),.A(g2459));
INVX1 NOT_4477 (.Y(g4377),.A(I7694));
INVX1 NOT_4478 (.Y(g4206),.A(I7435));
INVX1 NOT_4479 (.Y(I10651),.A(g6035));
INVX1 NOT_4480 (.Y(g3517),.A(I6702));
INVX1 NOT_4481 (.Y(g10575),.A(g10523));
INVX1 NOT_4482 (.Y(I14182),.A(g8788));
INVX1 NOT_4483 (.Y(I14672),.A(g9261));
INVX1 NOT_4484 (.Y(g7355),.A(I11713));
INVX1 NOT_4485 (.Y(g2045),.A(g1811));
INVX1 NOT_4486 (.Y(g7851),.A(g7479));
INVX1 NOT_4487 (.Y(I17549),.A(g11501));
INVX1 NOT_4488 (.Y(g3876),.A(I7061));
INVX1 NOT_4489 (.Y(g8131),.A(g8020));
INVX1 NOT_4490 (.Y(g10327),.A(I15771));
INVX1 NOT_4491 (.Y(g8331),.A(I13373));
INVX1 NOT_4492 (.Y(g2173),.A(I5120));
INVX1 NOT_4493 (.Y(I12120),.A(g7106));
INVX1 NOT_4494 (.Y(g2373),.A(g471));
INVX1 NOT_4495 (.Y(g4287),.A(I7546));
INVX1 NOT_4496 (.Y(I9276),.A(g5241));
INVX1 NOT_4497 (.Y(g10537),.A(I16178));
INVX1 NOT_4498 (.Y(I10331),.A(g6198));
INVX1 NOT_4499 (.Y(g7964),.A(g7651));
INVX1 NOT_4500 (.Y(g8635),.A(I13918));
INVX1 NOT_4501 (.Y(g6751),.A(I10762));
INVX1 NOT_4502 (.Y(I12562),.A(g7377));
INVX1 NOT_4503 (.Y(I8011),.A(g3820));
INVX1 NOT_4504 (.Y(I11947),.A(g6905));
INVX1 NOT_4505 (.Y(g8105),.A(g7992));
INVX1 NOT_4506 (.Y(g2169),.A(g42));
INVX1 NOT_4507 (.Y(I5395),.A(g892));
INVX1 NOT_4508 (.Y(I14449),.A(g8973));
INVX1 NOT_4509 (.Y(g10283),.A(g10166));
INVX1 NOT_4510 (.Y(g2369),.A(g617));
INVX1 NOT_4511 (.Y(I5913),.A(g2169));
INVX1 NOT_4512 (.Y(I11106),.A(g6667));
INVX1 NOT_4513 (.Y(g8487),.A(g8350));
INVX1 NOT_4514 (.Y(g2602),.A(I5707));
INVX1 NOT_4515 (.Y(I11605),.A(g6834));
INVX1 NOT_4516 (.Y(g4199),.A(I7414));
INVX1 NOT_4517 (.Y(g6585),.A(I10541));
INVX1 NOT_4518 (.Y(g2007),.A(g936));
INVX1 NOT_4519 (.Y(g5773),.A(I9359));
INVX1 NOT_4520 (.Y(g10492),.A(I16111));
INVX1 NOT_4521 (.Y(g4399),.A(g3638));
INVX1 NOT_4522 (.Y(g7463),.A(g6921));
INVX1 NOT_4523 (.Y(g2407),.A(g197));
INVX1 NOT_4524 (.Y(I6163),.A(g2547));
INVX1 NOT_4525 (.Y(g2920),.A(g2462));
INVX1 NOT_4526 (.Y(I14961),.A(g9769));
INVX1 NOT_4527 (.Y(g2578),.A(g1962));
INVX1 NOT_4528 (.Y(g2868),.A(I6010));
INVX1 NOT_4529 (.Y(g3214),.A(I6391));
INVX1 NOT_4530 (.Y(g4781),.A(I8147));
INVX1 NOT_4531 (.Y(g6041),.A(I9658));
INVX1 NOT_4532 (.Y(I6363),.A(g2459));
INVX1 NOT_4533 (.Y(I7202),.A(g2647));
INVX1 NOT_4534 (.Y(I15729),.A(g10254));
INVX1 NOT_4535 (.Y(I13812),.A(g8519));
INVX1 NOT_4536 (.Y(I9647),.A(g5148));
INVX1 NOT_4537 (.Y(g4898),.A(I8259));
INVX1 NOT_4538 (.Y(g6441),.A(g6151));
INVX1 NOT_4539 (.Y(I13463),.A(g8156));
INVX1 NOT_4540 (.Y(g9451),.A(I14642));
INVX1 NOT_4541 (.Y(g4900),.A(I8265));
INVX1 NOT_4542 (.Y(I6432),.A(g2350));
INVX1 NOT_4543 (.Y(g11501),.A(I17522));
INVX1 NOT_4544 (.Y(g3110),.A(g2482));
INVX1 NOT_4545 (.Y(g11577),.A(I17613));
INVX1 NOT_4546 (.Y(g7279),.A(g6382));
INVX1 NOT_4547 (.Y(g5836),.A(g5320));
INVX1 NOT_4548 (.Y(g4510),.A(I7909));
INVX1 NOT_4549 (.Y(g11439),.A(I17368));
INVX1 NOT_4550 (.Y(g3663),.A(I6832));
INVX1 NOT_4551 (.Y(I12427),.A(g7636));
INVX1 NOT_4552 (.Y(g10091),.A(I15320));
INVX1 NOT_4553 (.Y(g9346),.A(I14543));
INVX1 NOT_4554 (.Y(I12366),.A(g7134));
INVX1 NOT_4555 (.Y(g2261),.A(g1713));
INVX1 NOT_4556 (.Y(g7619),.A(I12205));
INVX1 NOT_4557 (.Y(g7318),.A(I11602));
INVX1 NOT_4558 (.Y(g2793),.A(g2276));
INVX1 NOT_4559 (.Y(g4291),.A(g4013));
INVX1 NOT_4560 (.Y(g7872),.A(I12655));
INVX1 NOT_4561 (.Y(g11438),.A(I17365));
INVX1 NOT_4562 (.Y(g10174),.A(I15514));
INVX1 NOT_4563 (.Y(g10796),.A(I16500));
INVX1 NOT_4564 (.Y(I16664),.A(g10795));
INVX1 NOT_4565 (.Y(g9103),.A(g8892));
INVX1 NOT_4566 (.Y(I8080),.A(g3538));
INVX1 NOT_4567 (.Y(g2015),.A(g1107));
INVX1 NOT_4568 (.Y(g6368),.A(g5987));
INVX1 NOT_4569 (.Y(g8445),.A(I13633));
INVX1 NOT_4570 (.Y(I7776),.A(g3773));
INVX1 NOT_4571 (.Y(g7057),.A(I11252));
INVX1 NOT_4572 (.Y(g2227),.A(g95));
INVX1 NOT_4573 (.Y(g4344),.A(g3946));
INVX1 NOT_4574 (.Y(I5142),.A(g639));
INVX1 NOT_4575 (.Y(I7593),.A(g4142));
INVX1 NOT_4576 (.Y(I5248),.A(g1110));
INVX1 NOT_4577 (.Y(g7989),.A(I12805));
INVX1 NOT_4578 (.Y(I9224),.A(g5063));
INVX1 NOT_4579 (.Y(I15284),.A(g10034));
INVX1 NOT_4580 (.Y(g3762),.A(I6965));
INVX1 NOT_4581 (.Y(I12403),.A(g7611));
INVX1 NOT_4582 (.Y(I12547),.A(g7673));
INVX1 NOT_4583 (.Y(g4207),.A(I7438));
INVX1 NOT_4584 (.Y(g11083),.A(g10913));
INVX1 NOT_4585 (.Y(g11348),.A(g11276));
INVX1 NOT_4586 (.Y(g10390),.A(g10309));
INVX1 NOT_4587 (.Y(I16484),.A(g10770));
INVX1 NOT_4588 (.Y(g9732),.A(I14873));
INVX1 NOT_4589 (.Y(I5815),.A(g1994));
INVX1 NOT_4590 (.Y(I9120),.A(g5218));
INVX1 NOT_4591 (.Y(g11284),.A(g11208));
INVX1 NOT_4592 (.Y(I9320),.A(g5013));
INVX1 NOT_4593 (.Y(g2246),.A(g1810));
INVX1 NOT_4594 (.Y(g5822),.A(g5320));
INVX1 NOT_4595 (.Y(g4819),.A(g3354));
INVX1 NOT_4596 (.Y(g3877),.A(I7064));
INVX1 NOT_4597 (.Y(g9508),.A(g9271));
INVX1 NOT_4598 (.Y(I12226),.A(g7066));
INVX1 NOT_4599 (.Y(g8007),.A(I12843));
INVX1 NOT_4600 (.Y(I7264),.A(g3252));
INVX1 NOT_4601 (.Y(g11622),.A(I17684));
INVX1 NOT_4602 (.Y(g2203),.A(g677));
INVX1 NOT_4603 (.Y(g7686),.A(g7148));
INVX1 NOT_4604 (.Y(g10192),.A(I15554));
INVX1 NOT_4605 (.Y(I10620),.A(g5884));
INVX1 NOT_4606 (.Y(I5497),.A(g587));
INVX1 NOT_4607 (.Y(I6929),.A(g2846));
INVX1 NOT_4608 (.Y(I12481),.A(g7570));
INVX1 NOT_4609 (.Y(I13421),.A(g8200));
INVX1 NOT_4610 (.Y(I16200),.A(g10494));
INVX1 NOT_4611 (.Y(g8868),.A(I14176));
INVX1 NOT_4612 (.Y(I5960),.A(g2239));
INVX1 NOT_4613 (.Y(I7360),.A(g4081));
INVX1 NOT_4614 (.Y(I14097),.A(g8773));
INVX1 NOT_4615 (.Y(I9617),.A(g5405));
INVX1 NOT_4616 (.Y(g6856),.A(I10924));
INVX1 NOT_4617 (.Y(g6411),.A(g6135));
INVX1 NOT_4618 (.Y(g6734),.A(I10733));
INVX1 NOT_4619 (.Y(I9789),.A(g5401));
INVX1 NOT_4620 (.Y(I10343),.A(g6003));
INVX1 NOT_4621 (.Y(g8535),.A(I13744));
INVX1 NOT_4622 (.Y(I7450),.A(g3704));
INVX1 NOT_4623 (.Y(I10971),.A(g6344));
INVX1 NOT_4624 (.Y(g7321),.A(I11611));
INVX1 NOT_4625 (.Y(g8582),.A(I13825));
INVX1 NOT_4626 (.Y(g7670),.A(I12289));
INVX1 NOT_4627 (.Y(I17261),.A(g11346));
INVX1 NOT_4628 (.Y(g4215),.A(I7462));
INVX1 NOT_4629 (.Y(I7996),.A(g3462));
INVX1 NOT_4630 (.Y(g11653),.A(I17761));
INVX1 NOT_4631 (.Y(g2502),.A(I5579));
INVX1 NOT_4632 (.Y(g4886),.A(I8231));
INVX1 NOT_4633 (.Y(g4951),.A(I8320));
INVX1 NOT_4634 (.Y(I16799),.A(g11017));
INVX1 NOT_4635 (.Y(g7232),.A(I11472));
INVX1 NOT_4636 (.Y(I12490),.A(g7637));
INVX1 NOT_4637 (.Y(g10553),.A(I16220));
INVX1 NOT_4638 (.Y(g8015),.A(I12857));
INVX1 NOT_4639 (.Y(I15415),.A(g10075));
INVX1 NOT_4640 (.Y(g5895),.A(g5361));
INVX1 NOT_4641 (.Y(g7938),.A(g7403));
INVX1 NOT_4642 (.Y(I8126),.A(g3662));
INVX1 NOT_4643 (.Y(g7813),.A(I12604));
INVX1 NOT_4644 (.Y(I5979),.A(g2543));
INVX1 NOT_4645 (.Y(g4314),.A(g4013));
INVX1 NOT_4646 (.Y(I5218),.A(g1104));
INVX1 NOT_4647 (.Y(g5062),.A(g4840));
INVX1 NOT_4648 (.Y(I13788),.A(g8517));
INVX1 NOT_4649 (.Y(g9347),.A(I14546));
INVX1 NOT_4650 (.Y(I12376),.A(g7195));
INVX1 NOT_4651 (.Y(g10326),.A(I15768));
INVX1 NOT_4652 (.Y(g5620),.A(g4417));
INVX1 NOT_4653 (.Y(g7909),.A(g7664));
INVX1 NOT_4654 (.Y(g2689),.A(g2038));
INVX1 NOT_4655 (.Y(I12103),.A(g6859));
INVX1 NOT_4656 (.Y(I11829),.A(g7213));
INVX1 NOT_4657 (.Y(g6863),.A(g6740));
INVX1 NOT_4658 (.Y(I16184),.A(g10484));
INVX1 NOT_4659 (.Y(I16805),.A(g10904));
INVX1 NOT_4660 (.Y(g10536),.A(I16175));
INVX1 NOT_4661 (.Y(g8664),.A(I13949));
INVX1 NOT_4662 (.Y(g10040),.A(I15247));
INVX1 NOT_4663 (.Y(I10412),.A(g5821));
INVX1 NOT_4664 (.Y(I12354),.A(g7143));
INVX1 NOT_4665 (.Y(g2216),.A(g41));
INVX1 NOT_4666 (.Y(g9533),.A(I14684));
INVX1 NOT_4667 (.Y(g6713),.A(I10698));
INVX1 NOT_4668 (.Y(I14412),.A(g8939));
INVX1 NOT_4669 (.Y(g7519),.A(g6956));
INVX1 NOT_4670 (.Y(I13828),.A(g8488));
INVX1 NOT_4671 (.Y(g10904),.A(I16664));
INVX1 NOT_4672 (.Y(g2028),.A(g1703));
INVX1 NOT_4673 (.Y(I14133),.A(g8772));
INVX1 NOT_4674 (.Y(g10252),.A(g10137));
INVX1 NOT_4675 (.Y(g8721),.A(g8582));
INVX1 NOT_4676 (.Y(g6569),.A(I10499));
INVX1 NOT_4677 (.Y(g10621),.A(I16298));
INVX1 NOT_4678 (.Y(g7606),.A(I12168));
INVX1 NOT_4679 (.Y(I6894),.A(g2813));
INVX1 NOT_4680 (.Y(I13344),.A(g8121));
INVX1 NOT_4681 (.Y(I10228),.A(g6113));
INVX1 NOT_4682 (.Y(g2247),.A(I5258));
INVX1 NOT_4683 (.Y(I14228),.A(g8797));
INVX1 NOT_4684 (.Y(g4336),.A(g4130));
INVX1 NOT_4685 (.Y(g3394),.A(I6598));
INVX1 NOT_4686 (.Y(I5830),.A(g2067));
INVX1 NOT_4687 (.Y(g2564),.A(g1814));
INVX1 NOT_4688 (.Y(g7687),.A(I12318));
INVX1 NOT_4689 (.Y(g4768),.A(I8126));
INVX1 NOT_4690 (.Y(g11576),.A(I17610));
INVX1 NOT_4691 (.Y(I10716),.A(g6093));
INVX1 NOT_4692 (.Y(I13682),.A(g8310));
INVX1 NOT_4693 (.Y(g3731),.A(I6911));
INVX1 NOT_4694 (.Y(I15554),.A(g10088));
INVX1 NOT_4695 (.Y(g2826),.A(g2163));
INVX1 NOT_4696 (.Y(I6661),.A(g2752));
INVX1 NOT_4697 (.Y(g6688),.A(I10655));
INVX1 NOT_4698 (.Y(I11173),.A(g6500));
INVX1 NOT_4699 (.Y(g10183),.A(g10042));
INVX1 NOT_4700 (.Y(g6857),.A(I10927));
INVX1 NOT_4701 (.Y(g5192),.A(g4640));
INVX1 NOT_4702 (.Y(g5085),.A(g4377));
INVX1 NOT_4703 (.Y(I5221),.A(g1407));
INVX1 NOT_4704 (.Y(g9820),.A(I14961));
INVX1 NOT_4705 (.Y(g4943),.A(I8311));
INVX1 NOT_4706 (.Y(I12190),.A(g7268));
INVX1 NOT_4707 (.Y(I7674),.A(g3352));
INVX1 NOT_4708 (.Y(g11200),.A(g11112));
INVX1 NOT_4709 (.Y(g10062),.A(I15284));
INVX1 NOT_4710 (.Y(g3705),.A(g3113));
INVX1 NOT_4711 (.Y(I16214),.A(g10500));
INVX1 NOT_4712 (.Y(I17271),.A(g11388));
INVX1 NOT_4713 (.Y(I12520),.A(g7415));
INVX1 NOT_4714 (.Y(g2638),.A(I5751));
INVX1 NOT_4715 (.Y(g4065),.A(g2794));
INVX1 NOT_4716 (.Y(I8161),.A(g3637));
INVX1 NOT_4717 (.Y(g4887),.A(I8234));
INVX1 NOT_4718 (.Y(g4228),.A(g3914));
INVX1 NOT_4719 (.Y(g4322),.A(I7593));
INVX1 NOT_4720 (.Y(g7570),.A(I12032));
INVX1 NOT_4721 (.Y(g2108),.A(I4992));
INVX1 NOT_4722 (.Y(g5941),.A(I9571));
INVX1 NOT_4723 (.Y(I14379),.A(g8961));
INVX1 NOT_4724 (.Y(g2609),.A(I5728));
INVX1 NOT_4725 (.Y(g4934),.A(g4243));
INVX1 NOT_4726 (.Y(g7341),.A(I11671));
INVX1 NOT_4727 (.Y(I11029),.A(g6485));
INVX1 NOT_4728 (.Y(g10851),.A(I16553));
INVX1 NOT_4729 (.Y(g10872),.A(I16586));
INVX1 NOT_4730 (.Y(g11052),.A(I16817));
INVX1 NOT_4731 (.Y(I5932),.A(g2539));
INVX1 NOT_4732 (.Y(I10958),.A(g6559));
INVX1 NOT_4733 (.Y(g6400),.A(I10308));
INVX1 NOT_4734 (.Y(I14112),.A(g8777));
INVX1 NOT_4735 (.Y(I10378),.A(g6244));
INVX1 NOT_4736 (.Y(g7525),.A(I11921));
INVX1 NOT_4737 (.Y(I7680),.A(g3736));
INVX1 NOT_4738 (.Y(I14958),.A(g9767));
INVX1 NOT_4739 (.Y(g2883),.A(I6037));
INVX1 NOT_4740 (.Y(g8671),.A(I13956));
INVX1 NOT_4741 (.Y(I6484),.A(g2073));
INVX1 NOT_4742 (.Y(I6439),.A(g2352));
INVX1 NOT_4743 (.Y(I9915),.A(g5304));
INVX1 NOT_4744 (.Y(g3254),.A(g2322));
INVX1 NOT_4745 (.Y(g9775),.A(g9474));
INVX1 NOT_4746 (.Y(I17736),.A(g11640));
INVX1 NOT_4747 (.Y(I15798),.A(g10281));
INVX1 NOT_4748 (.Y(g3814),.A(g3228));
INVX1 NOT_4749 (.Y(g5708),.A(I9253));
INVX1 NOT_4750 (.Y(I10096),.A(g5794));
INVX1 NOT_4751 (.Y(g2217),.A(I5192));
INVX1 NOT_4752 (.Y(g2758),.A(I5840));
INVX1 NOT_4753 (.Y(g5520),.A(I8943));
INVX1 NOT_4754 (.Y(I14944),.A(g9454));
INVX1 NOT_4755 (.Y(I17198),.A(g11319));
INVX1 NOT_4756 (.Y(I15184),.A(g9974));
INVX1 NOT_4757 (.Y(g4096),.A(I7236));
INVX1 NOT_4758 (.Y(g8564),.A(I13785));
INVX1 NOT_4759 (.Y(g3038),.A(g1982));
INVX1 NOT_4760 (.Y(g4496),.A(I7889));
INVX1 NOT_4761 (.Y(I8303),.A(g4784));
INVX1 NOT_4762 (.Y(g11184),.A(I16953));
INVX1 NOT_4763 (.Y(g5252),.A(g4640));
INVX1 NOT_4764 (.Y(g7607),.A(I12171));
INVX1 NOT_4765 (.Y(I17528),.A(g11487));
INVX1 NOT_4766 (.Y(I6702),.A(g2801));
INVX1 NOT_4767 (.Y(g3773),.A(I6996));
INVX1 NOT_4768 (.Y(g5812),.A(g5320));
INVX1 NOT_4769 (.Y(g3009),.A(g2135));
INVX1 NOT_4770 (.Y(I14681),.A(g9110));
INVX1 NOT_4771 (.Y(g2165),.A(I5098));
INVX1 NOT_4772 (.Y(g6183),.A(g5320));
INVX1 NOT_4773 (.Y(g2571),.A(g1822));
INVX1 NOT_4774 (.Y(g7659),.A(I12274));
INVX1 NOT_4775 (.Y(g2861),.A(I6001));
INVX1 NOT_4776 (.Y(g7358),.A(I11722));
INVX1 NOT_4777 (.Y(g4195),.A(I7402));
INVX1 NOT_4778 (.Y(g5176),.A(g4682));
INVX1 NOT_4779 (.Y(g6220),.A(g5446));
INVX1 NOT_4780 (.Y(I5716),.A(g2068));
INVX1 NOT_4781 (.Y(g10574),.A(I16239));
INVX1 NOT_4782 (.Y(I17764),.A(g11651));
INVX1 NOT_4783 (.Y(I5149),.A(g1453));
INVX1 NOT_4784 (.Y(g4395),.A(I7732));
INVX1 NOT_4785 (.Y(g10047),.A(I15266));
INVX1 NOT_4786 (.Y(g4337),.A(g4144));
INVX1 NOT_4787 (.Y(g4913),.A(I8285));
INVX1 NOT_4788 (.Y(I17365),.A(g11380));
INVX1 NOT_4789 (.Y(I14802),.A(g9666));
INVX1 NOT_4790 (.Y(g10205),.A(g10176));
INVX1 NOT_4791 (.Y(g2055),.A(g1950));
INVX1 NOT_4792 (.Y(g3769),.A(I6982));
INVX1 NOT_4793 (.Y(g10912),.A(I16688));
INVX1 NOT_4794 (.Y(g10311),.A(g10242));
INVX1 NOT_4795 (.Y(g2455),.A(g826));
INVX1 NOT_4796 (.Y(g9739),.A(I14884));
INVX1 NOT_4797 (.Y(g2827),.A(g2164));
INVX1 NOT_4798 (.Y(I6952),.A(g2867));
INVX1 NOT_4799 (.Y(I14793),.A(g9269));
INVX1 NOT_4800 (.Y(g3212),.A(I6385));
INVX1 NOT_4801 (.Y(I9402),.A(g5107));
INVX1 NOT_4802 (.Y(I12339),.A(g7054));
INVX1 NOT_4803 (.Y(I8240),.A(g4380));
INVX1 NOT_4804 (.Y(g1975),.A(g622));
INVX1 NOT_4805 (.Y(I5198),.A(g143));
INVX1 NOT_4806 (.Y(I12296),.A(g7236));
INVX1 NOT_4807 (.Y(g7311),.A(I11581));
INVX1 NOT_4808 (.Y(g2774),.A(g2276));
INVX1 NOT_4809 (.Y(I6616),.A(g3186));
INVX1 NOT_4810 (.Y(g3967),.A(g3247));
INVX1 NOT_4811 (.Y(I17161),.A(g11314));
INVX1 NOT_4812 (.Y(g6588),.A(I10546));
INVX1 NOT_4813 (.Y(I4935),.A(g585));
INVX1 NOT_4814 (.Y(I12644),.A(g7729));
INVX1 NOT_4815 (.Y(g2846),.A(I5970));
INVX1 NOT_4816 (.Y(I9762),.A(g5276));
INVX1 NOT_4817 (.Y(I10549),.A(g6184));
INVX1 NOT_4818 (.Y(g9079),.A(g8892));
INVX1 NOT_4819 (.Y(I13648),.A(g8376));
INVX1 NOT_4820 (.Y(g10051),.A(I15272));
INVX1 NOT_4821 (.Y(I14690),.A(g9150));
INVX1 NOT_4822 (.Y(g6161),.A(I9886));
INVX1 NOT_4823 (.Y(I14549),.A(g9262));
INVX1 NOT_4824 (.Y(g7615),.A(I12193));
INVX1 NOT_4825 (.Y(g6361),.A(g5867));
INVX1 NOT_4826 (.Y(g2196),.A(g91));
INVX1 NOT_4827 (.Y(g4266),.A(g3688));
INVX1 NOT_4828 (.Y(I7600),.A(g4159));
INVX1 NOT_4829 (.Y(g9668),.A(g9490));
INVX1 NOT_4830 (.Y(g2396),.A(g1389));
INVX1 NOT_4831 (.Y(g10592),.A(I16261));
INVX1 NOT_4832 (.Y(I15400),.A(g10069));
INVX1 NOT_4833 (.Y(g2803),.A(g2154));
INVX1 NOT_4834 (.Y(g5733),.A(I9287));
INVX1 NOT_4835 (.Y(I17225),.A(g11298));
DFFX1 DFF_82 (.CK(CK1), .D(g6812), .Q(g1098));
DFFX1 DFF_83 (.CK(CK1), .D(g8570), .Q(g932));
DFFX1 DFF_84 (.CK(CK1), .D(g5642), .Q(g126));
DFFX1 DFF_85 (.CK(CK1), .D(g8282), .Q(g1896));
DFFX1 DFF_86 (.CK(CK1), .D(g8435), .Q(g736));
DFFX1 DFF_87 (.CK(CK1), .D(g7807), .Q(g1019));
DFFX1 DFF_88 (.CK(CK1), .D(g7305), .Q(g1362));
DFFX1 DFF_89 (.CK(CK1), .D(g2639), .Q(g745));
DFFX1 DFF_90 (.CK(CK1), .D(g7332), .Q(g1419));
DFFX1 DFF_91 (.CK(CK1), .D(g7779), .Q(g58));
DFFX1 DFF_92 (.CK(CK1), .D(g11397), .Q(g32));
INVX1 NOT_4836 (.Y(g11400),.A(I17243));
INVX1 NOT_4837 (.Y(g6051),.A(I9680));
INVX1 NOT_4838 (.Y(I11770),.A(g7202));
INVX1 NOT_4839 (.Y(g5270),.A(g4367));
INVX1 NOT_4840 (.Y(g7374),.A(I11752));
INVX1 NOT_4841 (.Y(I11563),.A(g6819));
INVX1 NOT_4842 (.Y(I8116),.A(g3627));
INVX1 NOT_4843 (.Y(g6127),.A(I9826));
INVX1 NOT_4844 (.Y(g6451),.A(I10381));
INVX1 NOT_4845 (.Y(g8758),.A(I14055));
INVX1 NOT_4846 (.Y(g8066),.A(I12916));
INVX1 NOT_4847 (.Y(g8589),.A(I13834));
INVX1 NOT_4848 (.Y(I15329),.A(g9995));
INVX1 NOT_4849 (.Y(g7985),.A(I12799));
INVX1 NOT_4850 (.Y(I17258),.A(g11345));
INVX1 NOT_4851 (.Y(g4142),.A(I7288));
INVX1 NOT_4852 (.Y(g2509),.A(I5588));
INVX1 NOT_4853 (.Y(I16407),.A(g10696));
INVX1 NOT_4854 (.Y(I15539),.A(g10069));
INVX1 NOT_4855 (.Y(I6546),.A(g2987));
INVX1 NOT_4856 (.Y(g5073),.A(g4840));
INVX1 NOT_4857 (.Y(g10350),.A(I15814));
INVX1 NOT_4858 (.Y(g11207),.A(I16982));
INVX1 NOT_4859 (.Y(g1984),.A(g758));
INVX1 NOT_4860 (.Y(I10317),.A(g6003));
INVX1 NOT_4861 (.Y(g7284),.A(I11528));
INVX1 NOT_4862 (.Y(g11539),.A(g11519));
INVX1 NOT_4863 (.Y(g6146),.A(I9863));
INVX1 NOT_4864 (.Y(g10820),.A(I16528));
INVX1 NOT_4865 (.Y(g4081),.A(I7210));
INVX1 NOT_4866 (.Y(g7545),.A(I11967));
INVX1 NOT_4867 (.Y(g9356),.A(I14573));
INVX1 NOT_4868 (.Y(g8571),.A(I13806));
INVX1 NOT_4869 (.Y(I8147),.A(g3633));
INVX1 NOT_4870 (.Y(g2662),.A(g2014));
INVX1 NOT_4871 (.Y(g5124),.A(g4596));
INVX1 NOT_4872 (.Y(g2018),.A(g1336));
INVX1 NOT_4873 (.Y(g5980),.A(I9594));
INVX1 NOT_4874 (.Y(g2067),.A(g108));
INVX1 NOT_4875 (.Y(g7380),.A(g7279));
INVX1 NOT_4876 (.Y(g8448),.A(I13642));
INVX1 NOT_4877 (.Y(g6103),.A(I9766));
INVX1 NOT_4878 (.Y(I10129),.A(g5688));
INVX1 NOT_4879 (.Y(I9930),.A(g5317));
INVX1 NOT_4880 (.Y(I11767),.A(g7201));
INVX1 NOT_4881 (.Y(I11794),.A(g7188));
INVX1 NOT_4882 (.Y(g8711),.A(g8677));
INVX1 NOT_4883 (.Y(g7591),.A(I12103));
INVX1 NOT_4884 (.Y(g6303),.A(I10168));
INVX1 NOT_4885 (.Y(g2418),.A(I5497));
INVX1 NOT_4886 (.Y(I11845),.A(g6869));
INVX1 NOT_4887 (.Y(g5069),.A(g4368));
INVX1 NOT_4888 (.Y(I13794),.A(g8472));
INVX1 NOT_4889 (.Y(I10057),.A(g5741));
INVX1 NOT_4890 (.Y(g4726),.A(g3546));
INVX1 NOT_4891 (.Y(g2994),.A(g2057));
INVX1 NOT_4892 (.Y(g5469),.A(I8880));
INVX1 NOT_4893 (.Y(g7853),.A(I12652));
INVX1 NOT_4894 (.Y(g4354),.A(I7639));
INVX1 NOT_4895 (.Y(I5258),.A(g67));
INVX1 NOT_4896 (.Y(g7020),.A(I11159));
INVX1 NOT_4897 (.Y(I5818),.A(g2098));
INVX1 NOT_4898 (.Y(g8133),.A(I13002));
INVX1 NOT_4899 (.Y(g8333),.A(I13379));
INVX1 NOT_4900 (.Y(g7420),.A(I11804));
INVX1 NOT_4901 (.Y(I15241),.A(g10013));
INVX1 NOT_4902 (.Y(I11898),.A(g6896));
INVX1 NOT_4903 (.Y(g5177),.A(g4596));
INVX1 NOT_4904 (.Y(g6732),.A(I10729));
INVX1 NOT_4905 (.Y(I12867),.A(g7638));
INVX1 NOT_4906 (.Y(I17657),.A(g11598));
INVX1 NOT_4907 (.Y(I13633),.A(g8346));
INVX1 NOT_4908 (.Y(g11241),.A(g11112));
INVX1 NOT_4909 (.Y(I16206),.A(g10453));
INVX1 NOT_4910 (.Y(I10299),.A(g6243));
INVX1 NOT_4911 (.Y(g2256),.A(I5279));
INVX1 NOT_4912 (.Y(I11191),.A(g6514));
INVX1 NOT_4913 (.Y(I11719),.A(g7029));
INVX1 NOT_4914 (.Y(g7559),.A(I12009));
INVX1 NOT_4915 (.Y(I14323),.A(g8817));
INVX1 NOT_4916 (.Y(g10691),.A(I16360));
INVX1 NOT_4917 (.Y(g7794),.A(I12547));
INVX1 NOT_4918 (.Y(I7076),.A(g2985));
INVX1 NOT_4919 (.Y(I13191),.A(g8132));
INVX1 NOT_4920 (.Y(I14299),.A(g8810));
INVX1 NOT_4921 (.Y(I7889),.A(g3373));
INVX1 NOT_4922 (.Y(g8196),.A(I13125));
INVX1 NOT_4923 (.Y(g6944),.A(I11082));
INVX1 NOT_4924 (.Y(g8803),.A(I14130));
INVX1 NOT_4925 (.Y(I6277),.A(g1206));
INVX1 NOT_4926 (.Y(g6072),.A(g4977));
INVX1 NOT_4927 (.Y(I15771),.A(g10250));
INVX1 NOT_4928 (.Y(I9237),.A(g5205));
INVX1 NOT_4929 (.Y(I17337),.A(g11363));
INVX1 NOT_4930 (.Y(g2181),.A(I5142));
INVX1 NOT_4931 (.Y(g8538),.A(I13747));
INVX1 NOT_4932 (.Y(g2381),.A(g1368));
INVX1 NOT_4933 (.Y(g9432),.A(g9313));
INVX1 NOT_4934 (.Y(I15235),.A(g9968));
INVX1 NOT_4935 (.Y(I6789),.A(g2748));
INVX1 NOT_4949 (.Y(g2197),.A(g101));
INVX1 NOT_4950 (.Y(I7651),.A(g3332));
INVX1 NOT_4951 (.Y(g4312),.A(g4144));
INVX1 NOT_4952 (.Y(I8820),.A(g4473));
INVX1 NOT_4953 (.Y(I11440),.A(g6577));
INVX1 NOT_4954 (.Y(g10929),.A(g10827));
INVX1 NOT_4955 (.Y(I12496),.A(g7724));
INVX1 NOT_4956 (.Y(g2021),.A(g1341));
INVX1 NOT_4957 (.Y(I9194),.A(g5236));
INVX1 NOT_4958 (.Y(g7628),.A(I12226));
INVX1 NOT_4959 (.Y(I9394),.A(g5195));
INVX1 NOT_4960 (.Y(g6116),.A(I9801));
INVX1 NOT_4961 (.Y(g2421),.A(g1374));
INVX1 NOT_4962 (.Y(g7630),.A(I12232));
INVX1 NOT_4963 (.Y(g4001),.A(g3200));
INVX1 NOT_4964 (.Y(I12978),.A(g8040));
INVX1 NOT_4965 (.Y(I14232),.A(g8800));
INVX1 NOT_4966 (.Y(g10928),.A(g10827));
INVX1 NOT_4967 (.Y(g8067),.A(I12919));
INVX1 NOT_4968 (.Y(I9731),.A(g5255));
INVX1 NOT_4969 (.Y(g5898),.A(g5361));
INVX1 NOT_4970 (.Y(g8418),.A(I13568));
INVX1 NOT_4971 (.Y(g6434),.A(I10352));
INVX1 NOT_4972 (.Y(g4676),.A(g3354));
INVX1 NOT_4973 (.Y(g5900),.A(I9531));
INVX1 NOT_4974 (.Y(g6565),.A(g5790));
INVX1 NOT_4975 (.Y(I5821),.A(g2101));
INVX1 NOT_4976 (.Y(I6299),.A(g2242));
INVX1 NOT_4977 (.Y(I11926),.A(g6900));
INVX1 NOT_4978 (.Y(g8290),.A(I13224));
INVX1 NOT_4979 (.Y(I12986),.A(g8042));
INVX1 NOT_4980 (.Y(g4129),.A(I7280));
INVX1 NOT_4981 (.Y(g5797),.A(I9399));
INVX1 NOT_4982 (.Y(g4329),.A(g4144));
INVX1 NOT_4983 (.Y(I14697),.A(g9260));
INVX1 NOT_4984 (.Y(g4761),.A(g3440));
INVX1 NOT_4985 (.Y(g11515),.A(g11490));
INVX1 NOT_4986 (.Y(I7384),.A(g4082));
INVX1 NOT_4987 (.Y(I13612),.A(g8325));
INVX1 NOT_4988 (.Y(g5245),.A(g4369));
INVX1 NOT_4989 (.Y(I7339),.A(g4004));
INVX1 NOT_4990 (.Y(I13099),.A(g7927));
INVX1 NOT_4991 (.Y(I12384),.A(g7212));
INVX1 NOT_4992 (.Y(g8093),.A(I12948));
INVX1 NOT_4993 (.Y(I13388),.A(g8230));
INVX1 NOT_4994 (.Y(g6681),.A(g5830));
INVX1 NOT_4995 (.Y(I11701),.A(g7065));
INVX1 NOT_4996 (.Y(I11534),.A(g6917));
INVX1 NOT_4997 (.Y(g10787),.A(I16487));
INVX1 NOT_4998 (.Y(g5291),.A(g4384));
INVX1 NOT_4999 (.Y(g3392),.A(g3121));
INVX1 NOT_5000 (.Y(I11272),.A(g6546));
INVX1 NOT_5001 (.Y(g10282),.A(g10164));
INVX1 NOT_5002 (.Y(g7750),.A(I12415));
INVX1 NOT_5003 (.Y(g3485),.A(g2662));
INVX1 NOT_5004 (.Y(g2562),.A(g1383));
INVX1 NOT_5005 (.Y(g6697),.A(g5949));
INVX1 NOT_5006 (.Y(g5144),.A(g4682));
INVX1 NOT_5007 (.Y(g4592),.A(g3829));
INVX1 NOT_5008 (.Y(g6914),.A(I11024));
INVX1 NOT_5009 (.Y(I17444),.A(g11446));
INVX1 NOT_5010 (.Y(g5344),.A(I8811));
INVX1 NOT_5011 (.Y(g6210),.A(g5205));
INVX1 NOT_5012 (.Y(I12150),.A(g7074));
INVX1 NOT_5013 (.Y(g4746),.A(I8098));
INVX1 NOT_5014 (.Y(g8181),.A(I13096));
INVX1 NOT_5015 (.Y(g10827),.A(I16543));
INVX1 NOT_5016 (.Y(g6596),.A(I10566));
INVX1 NOT_5017 (.Y(I6738),.A(g3113));
INVX1 NOT_5018 (.Y(g4221),.A(g3914));
INVX1 NOT_5019 (.Y(g8381),.A(I13489));
INVX1 NOT_5020 (.Y(g2101),.A(I4951));
INVX1 NOT_5021 (.Y(g2817),.A(I5919));
INVX1 NOT_5022 (.Y(g3941),.A(g3015));
INVX1 NOT_5023 (.Y(g7040),.A(I11207));
INVX1 NOT_5024 (.Y(g6413),.A(I10325));
INVX1 NOT_5025 (.Y(I10831),.A(g6710));
INVX1 NOT_5026 (.Y(g7440),.A(I11836));
INVX1 NOT_5027 (.Y(g8197),.A(I13128));
INVX1 NOT_5028 (.Y(g8700),.A(g8574));
INVX1 NOT_5029 (.Y(I10445),.A(g5770));
INVX1 NOT_5030 (.Y(I7523),.A(g4095));
INVX1 NOT_5031 (.Y(I11140),.A(g6448));
INVX1 NOT_5032 (.Y(I12196),.A(g7272));
INVX1 NOT_5033 (.Y(g2605),.A(I5716));
INVX1 NOT_5034 (.Y(g11441),.A(I17374));
INVX1 NOT_5035 (.Y(I9150),.A(g5012));
INVX1 NOT_5036 (.Y(I10499),.A(g6149));
INVX1 NOT_5037 (.Y(g8421),.A(I13577));
INVX1 NOT_5038 (.Y(g7123),.A(I11360));
INVX1 NOT_5039 (.Y(g5088),.A(I8456));
INVX1 NOT_5040 (.Y(g11206),.A(I16979));
INVX1 NOT_5041 (.Y(g7323),.A(I11617));
INVX1 NOT_5042 (.Y(I14499),.A(g8889));
INVX1 NOT_5043 (.Y(I6907),.A(g2994));
INVX1 NOT_5044 (.Y(I12526),.A(g7648));
INVX1 NOT_5045 (.Y(g10803),.A(g10708));
INVX1 NOT_5046 (.Y(I7205),.A(g2632));
INVX1 NOT_5047 (.Y(I9773),.A(g4934));
INVX1 NOT_5048 (.Y(I15759),.A(g10267));
INVX1 NOT_5049 (.Y(I11061),.A(g6641));
INVX1 NOT_5050 (.Y(I15725),.A(g10251));
INVX1 NOT_5051 (.Y(g5701),.A(I9240));
INVX1 NOT_5052 (.Y(g3708),.A(I6867));
INVX1 NOT_5053 (.Y(g4953),.A(I8324));
INVX1 NOT_5054 (.Y(g2751),.A(I5821));
INVX1 NOT_5055 (.Y(g3520),.A(g2779));
INVX1 NOT_5056 (.Y(g8950),.A(I14303));
INVX1 NOT_5057 (.Y(I16500),.A(g10711));
INVX1 NOT_5058 (.Y(g3219),.A(I6395));
INVX1 NOT_5059 (.Y(I6517),.A(g3271));
INVX1 NOT_5060 (.Y(I6690),.A(g2743));
INVX1 NOT_5061 (.Y(I9409),.A(g5013));
INVX1 NOT_5062 (.Y(I15114),.A(g9875));
INVX1 NOT_5063 (.Y(I5427),.A(g913));
INVX1 NOT_5064 (.Y(g4468),.A(I7837));
INVX1 NOT_5065 (.Y(I15082),.A(g9719));
INVX1 NOT_5066 (.Y(g6117),.A(I9804));
INVX1 NOT_5067 (.Y(I14989),.A(g9813));
INVX1 NOT_5068 (.Y(I17158),.A(g11312));
INVX1 NOT_5069 (.Y(g3252),.A(I6414));
INVX1 NOT_5070 (.Y(g10881),.A(I16613));
INVX1 NOT_5071 (.Y(I7104),.A(g3186));
INVX1 NOT_5072 (.Y(g11435),.A(I17356));
INVX1 NOT_5073 (.Y(I6876),.A(g2956));
INVX1 NOT_5074 (.Y(I9769),.A(g5287));
INVX1 NOT_5075 (.Y(g11082),.A(I16859));
INVX1 NOT_5076 (.Y(g3812),.A(g3228));
INVX1 NOT_5077 (.Y(I7099),.A(g3228));
INVX1 NOT_5078 (.Y(I12457),.A(g7559));
INVX1 NOT_5079 (.Y(I10924),.A(g6736));
INVX1 NOT_5080 (.Y(g5886),.A(g5361));
INVX1 NOT_5081 (.Y(g11107),.A(g10974));
INVX1 NOT_5082 (.Y(I9836),.A(g5405));
INVX1 NOT_5083 (.Y(I14080),.A(g8714));
INVX1 NOT_5084 (.Y(g7351),.A(I11701));
INVX1 NOT_5085 (.Y(g2041),.A(g1791));
INVX1 NOT_5086 (.Y(g7648),.A(I12255));
INVX1 NOT_5087 (.Y(g7530),.A(I11926));
INVX1 NOT_5088 (.Y(I11360),.A(g6351));
INVX1 NOT_5089 (.Y(g8562),.A(I13779));
INVX1 NOT_5090 (.Y(I15744),.A(g10261));
INVX1 NOT_5091 (.Y(I13360),.A(g8126));
INVX1 NOT_5092 (.Y(I17353),.A(g11381));
INVX1 NOT_5093 (.Y(g3405),.A(g3144));
INVX1 NOT_5094 (.Y(g5114),.A(I8506));
INVX1 NOT_5095 (.Y(I5403),.A(g636));
INVX1 NOT_5096 (.Y(g9778),.A(g9474));
INVX1 NOT_5097 (.Y(g5314),.A(g4387));
INVX1 NOT_5098 (.Y(I11447),.A(g6431));
INVX1 NOT_5099 (.Y(g11345),.A(I17158));
INVX1 NOT_5100 (.Y(g9894),.A(I15085));
INVX1 NOT_5101 (.Y(g8723),.A(g8585));
INVX1 NOT_5102 (.Y(g4716),.A(g3546));
INVX1 NOT_5103 (.Y(I11162),.A(g6479));
INVX1 NOT_5104 (.Y(I16613),.A(g10794));
INVX1 NOT_5105 (.Y(g11399),.A(I17240));
INVX1 NOT_5106 (.Y(g3765),.A(g3120));
INVX1 NOT_5107 (.Y(I10753),.A(g5814));
INVX1 NOT_5108 (.Y(I10461),.A(g5849));
INVX1 NOT_5109 (.Y(I5391),.A(g1101));
INVX1 NOT_5110 (.Y(g3911),.A(g3015));
INVX1 NOT_5111 (.Y(I9229),.A(g4954));
INVX1 NOT_5112 (.Y(g7010),.A(I11155));
INVX1 NOT_5113 (.Y(g6581),.A(I10531));
INVX1 NOT_5114 (.Y(g10890),.A(I16632));
INVX1 NOT_5115 (.Y(g5650),.A(I9111));
INVX1 NOT_5116 (.Y(g7410),.A(I11790));
INVX1 NOT_5117 (.Y(g9782),.A(I14933));
INVX1 NOT_5118 (.Y(g11398),.A(I17237));
INVX1 NOT_5119 (.Y(I15804),.A(g10283));
INVX1 NOT_5120 (.Y(I16947),.A(g11080));
INVX1 NOT_5121 (.Y(I5695),.A(g575));
INVX1 NOT_5122 (.Y(g10249),.A(g10135));
INVX1 NOT_5123 (.Y(g2168),.A(I5111));
INVX1 NOT_5124 (.Y(g2669),.A(g2015));
INVX1 NOT_5125 (.Y(g6060),.A(I9695));
INVX1 NOT_5126 (.Y(I16273),.A(g10559));
INVX1 NOT_5127 (.Y(g2368),.A(I5445));
INVX1 NOT_5128 (.Y(I11629),.A(g6914));
INVX1 NOT_5129 (.Y(g11652),.A(I17758));
INVX1 NOT_5130 (.Y(I9822),.A(g5219));
INVX1 NOT_5131 (.Y(g9661),.A(I14786));
INVX1 NOT_5132 (.Y(g4198),.A(I7411));
INVX1 NOT_5133 (.Y(g4747),.A(g3586));
INVX1 NOT_5134 (.Y(I11472),.A(g6488));
INVX1 NOT_5135 (.Y(I10736),.A(g6104));
INVX1 NOT_5136 (.Y(g4398),.A(g3914));
INVX1 NOT_5137 (.Y(I13451),.A(g8152));
INVX1 NOT_5138 (.Y(g3733),.A(I6917));
INVX1 NOT_5139 (.Y(I7444),.A(g3683));
INVX1 NOT_5140 (.Y(g10248),.A(g10134));
INVX1 NOT_5141 (.Y(g2772),.A(g2508));
INVX1 NOT_5142 (.Y(I7269),.A(g2851));
INVX1 NOT_5143 (.Y(I15263),.A(g9995));
INVX1 NOT_5144 (.Y(I10198),.A(g6118));
INVX1 NOT_5145 (.Y(I12300),.A(g7240));
INVX1 NOT_5146 (.Y(g10552),.A(I16217));
INVX1 NOT_5147 (.Y(g8751),.A(g8632));
INVX1 NOT_5148 (.Y(I15332),.A(g10001));
INVX1 NOT_5149 (.Y(g10204),.A(g10174));
INVX1 NOT_5150 (.Y(g2743),.A(I5801));
INVX1 NOT_5151 (.Y(g4241),.A(g3664));
INVX1 NOT_5152 (.Y(g2890),.A(I6052));
INVX1 NOT_5153 (.Y(g5768),.A(I9352));
INVX1 NOT_5154 (.Y(I10843),.A(g6723));
INVX1 NOT_5155 (.Y(g8585),.A(I13828));
INVX1 NOT_5156 (.Y(I5858),.A(g2529));
INVX1 NOT_5157 (.Y(g5594),.A(I9016));
INVX1 NOT_5158 (.Y(I14528),.A(g9270));
INVX1 NOT_5159 (.Y(g3473),.A(I6676));
INVX1 NOT_5160 (.Y(g7278),.A(I11524));
INVX1 NOT_5161 (.Y(I14330),.A(g8819));
INVX1 NOT_5162 (.Y(g9526),.A(g9256));
INVX1 NOT_5163 (.Y(I4938),.A(g261));
INVX1 NOT_5164 (.Y(I8250),.A(g4589));
INVX1 NOT_5165 (.Y(I11071),.A(g6656));
INVX1 NOT_5166 (.Y(I15406),.A(g10065));
INVX1 NOT_5167 (.Y(I15962),.A(g10405));
INVX1 NOT_5168 (.Y(g2011),.A(g976));
INVX1 NOT_5169 (.Y(g6995),.A(g6482));
INVX1 NOT_5170 (.Y(g7618),.A(I12202));
INVX1 NOT_5171 (.Y(g3980),.A(g3121));
INVX1 NOT_5172 (.Y(g8441),.A(I13621));
INVX1 NOT_5173 (.Y(g11406),.A(I17261));
INVX1 NOT_5174 (.Y(g5943),.A(I9581));
INVX1 NOT_5175 (.Y(g7343),.A(I11677));
INVX1 NOT_5176 (.Y(g2411),.A(I5494));
INVX1 NOT_5177 (.Y(I10132),.A(g5696));
INVX1 NOT_5178 (.Y(g10786),.A(I16484));
INVX1 NOT_5179 (.Y(g3069),.A(I6277));
INVX1 NOT_5180 (.Y(I13776),.A(g8513));
INVX1 NOT_5181 (.Y(I13785),.A(g8516));
INVX1 NOT_5182 (.Y(g1982),.A(g736));
INVX1 NOT_5183 (.Y(g4524),.A(g3946));
INVX1 NOT_5184 (.Y(g6294),.A(I10141));
INVX1 NOT_5185 (.Y(I15500),.A(g10051));
INVX1 NOT_5186 (.Y(I5251),.A(g1424));
INVX1 NOT_5187 (.Y(I6590),.A(g3186));
INVX1 NOT_5188 (.Y(g3540),.A(g3307));
INVX1 NOT_5189 (.Y(I7729),.A(g3757));
INVX1 NOT_5190 (.Y(g5887),.A(I9510));
INVX1 NOT_5191 (.Y(g10356),.A(I15832));
INVX1 NOT_5192 (.Y(I5047),.A(g1185));
INVX1 NOT_5193 (.Y(g5122),.A(g4682));
INVX1 NOT_5194 (.Y(g11500),.A(I17519));
INVX1 NOT_5195 (.Y(g6190),.A(g5426));
INVX1 NOT_5196 (.Y(g2074),.A(g1377));
INVX1 NOT_5197 (.Y(g4319),.A(g4144));
INVX1 NOT_5198 (.Y(g7693),.A(I12326));
INVX1 NOT_5199 (.Y(g11049),.A(I16808));
INVX1 NOT_5200 (.Y(I11950),.A(g6906));
INVX1 NOT_5201 (.Y(I16514),.A(g10717));
INVX1 NOT_5202 (.Y(g10826),.A(I16540));
INVX1 NOT_5203 (.Y(I9062),.A(g4759));
INVX1 NOT_5204 (.Y(g7334),.A(I11650));
INVX1 NOT_5205 (.Y(g10380),.A(I15864));
INVX1 NOT_5206 (.Y(g3206),.A(g2055));
INVX1 NOT_5207 (.Y(I13825),.A(g8488));
INVX1 NOT_5208 (.Y(I13370),.A(g8128));
INVX1 NOT_5209 (.Y(I9620),.A(g5189));
INVX1 NOT_5210 (.Y(g4258),.A(I7509));
INVX1 NOT_5211 (.Y(I16507),.A(g10712));
INVX1 NOT_5212 (.Y(g4352),.A(I7633));
INVX1 NOT_5213 (.Y(I11858),.A(g6888));
INVX1 NOT_5214 (.Y(g11048),.A(I16805));
INVX1 NOT_5215 (.Y(g4577),.A(I7984));
INVX1 NOT_5216 (.Y(g4867),.A(I8204));
INVX1 NOT_5217 (.Y(I14709),.A(g9267));
INVX1 NOT_5218 (.Y(g5033),.A(I8406));
INVX1 NOT_5219 (.Y(g10233),.A(g10187));
INVX1 NOT_5220 (.Y(g6156),.A(g5426));
INVX1 NOT_5221 (.Y(g4717),.A(g3829));
INVX1 NOT_5222 (.Y(I7014),.A(g2919));
INVX1 NOT_5223 (.Y(I12511),.A(g7733));
INVX1 NOT_5224 (.Y(g10182),.A(I15530));
INVX1 NOT_5225 (.Y(g7555),.A(I11989));
INVX1 NOT_5226 (.Y(g7804),.A(I12577));
INVX1 NOT_5227 (.Y(I7414),.A(g4156));
INVX1 NOT_5228 (.Y(I10087),.A(g5753));
INVX1 NOT_5229 (.Y(g9919),.A(I15114));
INVX1 NOT_5230 (.Y(g2080),.A(I4894));
INVX1 NOT_5231 (.Y(I7946),.A(g3417));
INVX1 NOT_5232 (.Y(I10258),.A(g6134));
INVX1 NOT_5233 (.Y(I14087),.A(g8770));
INVX1 NOT_5234 (.Y(g7792),.A(I12541));
INVX1 NOT_5235 (.Y(g2480),.A(I5561));
INVX1 NOT_5236 (.Y(I11367),.A(g6392));
INVX1 NOT_5237 (.Y(I11394),.A(g6621));
INVX1 NOT_5238 (.Y(g5096),.A(g4840));
INVX1 NOT_5239 (.Y(g6942),.A(I11076));
INVX1 NOT_5240 (.Y(g8890),.A(I14236));
INVX1 NOT_5241 (.Y(g2713),.A(g2042));
INVX1 NOT_5242 (.Y(I13367),.A(g8221));
INVX1 NOT_5243 (.Y(I13394),.A(g8137));
INVX1 NOT_5244 (.Y(g4211),.A(I7450));
INVX1 NOT_5245 (.Y(g4186),.A(I7375));
INVX1 NOT_5246 (.Y(g6704),.A(g5949));
INVX1 NOT_5247 (.Y(I17687),.A(g11610));
INVX1 NOT_5248 (.Y(g4386),.A(I7713));
INVX1 NOT_5249 (.Y(g10932),.A(g10827));
INVX1 NOT_5250 (.Y(I8929),.A(g4582));
INVX1 NOT_5251 (.Y(g5845),.A(g5320));
INVX1 NOT_5252 (.Y(g4975),.A(I8351));
INVX1 NOT_5253 (.Y(g2569),.A(I5695));
INVX1 NOT_5254 (.Y(I7513),.A(g4144));
INVX1 NOT_5255 (.Y(g8011),.A(I12853));
INVX1 NOT_5256 (.Y(I17752),.A(g11645));
INVX1 NOT_5257 (.Y(g5195),.A(g4453));
INVX1 NOT_5258 (.Y(g5395),.A(I8831));
INVX1 NOT_5259 (.Y(g5891),.A(g5361));
INVX1 NOT_5260 (.Y(I9842),.A(g5405));
INVX1 NOT_5261 (.Y(I17374),.A(g11411));
INVX1 NOT_5262 (.Y(g7113),.A(I11348));
INVX1 NOT_5263 (.Y(g11106),.A(g10974));
INVX1 NOT_5264 (.Y(g7313),.A(I11587));
INVX1 NOT_5265 (.Y(I11420),.A(g6417));
INVX1 NOT_5266 (.Y(g4426),.A(g3914));
INVX1 NOT_5267 (.Y(g10897),.A(g10827));
INVX1 NOT_5268 (.Y(I12916),.A(g7849));
INVX1 NOT_5269 (.Y(I10069),.A(g5787));
INVX1 NOT_5270 (.Y(g6954),.A(I11100));
INVX1 NOT_5271 (.Y(g6250),.A(I10009));
INVX1 NOT_5272 (.Y(g4170),.A(g3328));
INVX1 NOT_5273 (.Y(g6810),.A(I10840));
INVX1 NOT_5274 (.Y(g4614),.A(g3829));
INVX1 NOT_5275 (.Y(g9527),.A(I14668));
INVX1 NOT_5276 (.Y(g4370),.A(I7671));
INVX1 NOT_5277 (.Y(I12550),.A(g7675));
INVX1 NOT_5278 (.Y(I7378),.A(g4067));
INVX1 NOT_5279 (.Y(I10810),.A(g6539));
INVX1 NOT_5280 (.Y(I11318),.A(g6488));
INVX1 NOT_5281 (.Y(g4125),.A(I7272));
INVX1 NOT_5282 (.Y(I15371),.A(g9990));
INVX1 NOT_5283 (.Y(g6432),.A(g6146));
INVX1 NOT_5284 (.Y(g7908),.A(g7454));
INVX1 NOT_5285 (.Y(I13227),.A(g8264));
INVX1 NOT_5286 (.Y(g6053),.A(I9684));
INVX1 NOT_5287 (.Y(I14955),.A(g9765));
INVX1 NOT_5288 (.Y(I17669),.A(g11604));
INVX1 NOT_5289 (.Y(g8992),.A(I14397));
INVX1 NOT_5290 (.Y(g9764),.A(g9432));
INVX1 NOT_5291 (.Y(I16920),.A(g11084));
INVX1 NOT_5292 (.Y(g11033),.A(I16760));
INVX1 NOT_5293 (.Y(g3291),.A(g2161));
INVX1 NOT_5294 (.Y(I12307),.A(g7245));
INVX1 NOT_5295 (.Y(I5935),.A(g2174));
INVX1 NOT_5296 (.Y(I6844),.A(g2915));
INVX1 NOT_5297 (.Y(g6453),.A(g5817));
INVX1 NOT_5298 (.Y(I9854),.A(g5557));
INVX1 NOT_5299 (.Y(I14970),.A(g9732));
INVX1 NOT_5300 (.Y(g4280),.A(g4013));
INVX1 NOT_5301 (.Y(I7182),.A(g2645));
INVX1 NOT_5302 (.Y(I7288),.A(g2873));
INVX1 NOT_5303 (.Y(g4939),.A(I8303));
INVX1 NOT_5304 (.Y(I11540),.A(g6877));
INVX1 NOT_5305 (.Y(I5982),.A(g2510));
INVX1 NOT_5306 (.Y(g3144),.A(g2462));
INVX1 NOT_5307 (.Y(I11058),.A(g6641));
INVX1 NOT_5308 (.Y(I15795),.A(g10280));
INVX1 NOT_5309 (.Y(g3344),.A(I6528));
INVX1 NOT_5310 (.Y(I16121),.A(g10396));
INVX1 NOT_5311 (.Y(g6568),.A(g5797));
INVX1 NOT_5312 (.Y(I10171),.A(g5992));
INVX1 NOT_5313 (.Y(g4083),.A(I7216));
INVX1 NOT_5314 (.Y(g8080),.A(I12942));
INVX1 NOT_5315 (.Y(I4879),.A(g256));
INVX1 NOT_5316 (.Y(g4544),.A(g3880));
INVX1 NOT_5317 (.Y(g3207),.A(g2439));
INVX1 NOT_5318 (.Y(g8573),.A(I13812));
INVX1 NOT_5319 (.Y(I7916),.A(g3664));
INVX1 NOT_5320 (.Y(I7022),.A(g2941));
INVX1 NOT_5321 (.Y(I13203),.A(g8196));
INVX1 NOT_5322 (.Y(g8480),.A(I13682));
INVX1 NOT_5323 (.Y(g7776),.A(I12493));
INVX1 NOT_5324 (.Y(g2000),.A(g810));
INVX1 NOT_5325 (.Y(I7749),.A(g3764));
INVX1 NOT_5326 (.Y(I6557),.A(g3086));
INVX1 NOT_5327 (.Y(g8713),.A(g8684));
INVX1 NOT_5328 (.Y(I17525),.A(g11486));
INVX1 NOT_5329 (.Y(g2126),.A(g12));
INVX1 NOT_5330 (.Y(g4636),.A(I8036));
INVX1 NOT_5331 (.Y(I15514),.A(g10122));
INVX1 NOT_5332 (.Y(I17424),.A(g11424));
INVX1 NOT_5333 (.Y(g3694),.A(I6851));
INVX1 NOT_5334 (.Y(g6157),.A(I9880));
INVX1 NOT_5335 (.Y(I6071),.A(g2269));
INVX1 NOT_5336 (.Y(I14967),.A(g9763));
INVX1 NOT_5337 (.Y(I12773),.A(g7581));
INVX1 NOT_5338 (.Y(I16682),.A(g10799));
INVX1 NOT_5339 (.Y(I17558),.A(g11504));
INVX1 NOT_5340 (.Y(I15507),.A(g10047));
INVX1 NOT_5341 (.Y(g5081),.A(I8449));
INVX1 NOT_5342 (.Y(I12942),.A(g7982));
INVX1 NOT_5343 (.Y(g3088),.A(I6294));
INVX1 NOT_5344 (.Y(g5815),.A(I9421));
INVX1 NOT_5345 (.Y(g8569),.A(I13800));
INVX1 NOT_5346 (.Y(g4306),.A(g3586));
INVX1 NOT_5347 (.Y(g7965),.A(I12759));
INVX1 NOT_5348 (.Y(I12268),.A(g7107));
INVX1 NOT_5349 (.Y(g5481),.A(I8900));
INVX1 NOT_5350 (.Y(g11507),.A(I17540));
INVX1 NOT_5351 (.Y(I12156),.A(g6878));
INVX1 NOT_5352 (.Y(g4790),.A(g3337));
INVX1 NOT_5353 (.Y(I12655),.A(g7402));
INVX1 NOT_5354 (.Y(g5692),.A(I9221));
INVX1 NOT_5355 (.Y(I15421),.A(g10083));
INVX1 NOT_5356 (.Y(g1964),.A(g114));
INVX1 NOT_5357 (.Y(g10387),.A(g10357));
INVX1 NOT_5358 (.Y(g97),.A(I4780));
INVX1 NOT_5359 (.Y(g7264),.A(I11501));
INVX1 NOT_5360 (.Y(I12180),.A(g7263));
INVX1 NOT_5361 (.Y(g10620),.A(I16295));
INVX1 NOT_5362 (.Y(g4187),.A(I7378));
INVX1 NOT_5363 (.Y(g4061),.A(I7182));
INVX1 NOT_5364 (.Y(g10148),.A(g10121));
INVX1 NOT_5365 (.Y(g11421),.A(I17318));
INVX1 NOT_5366 (.Y(g4387),.A(I7716));
INVX1 NOT_5367 (.Y(g4461),.A(g3829));
INVX1 NOT_5368 (.Y(I6955),.A(g2871));
INVX1 NOT_5369 (.Y(g7360),.A(I11728));
INVX1 NOT_5370 (.Y(g11163),.A(I16920));
INVX1 NOT_5371 (.Y(g10104),.A(I15338));
INVX1 NOT_5372 (.Y(I11146),.A(g6439));
INVX1 NOT_5373 (.Y(g4756),.A(g3440));
INVX1 NOT_5374 (.Y(I17713),.A(g11621));
INVX1 NOT_5375 (.Y(I13738),.A(g8295));
INVX1 NOT_5376 (.Y(I13645),.A(g8379));
INVX1 NOT_5377 (.Y(g8688),.A(g8507));
INVX1 NOT_5378 (.Y(I12335),.A(g7133));
INVX1 NOT_5379 (.Y(g7521),.A(I11901));
INVX1 NOT_5380 (.Y(g10343),.A(I15795));
INVX1 NOT_5381 (.Y(I14010),.A(g8642));
INVX1 NOT_5382 (.Y(I14918),.A(g9535));
INVX1 NOT_5383 (.Y(g8976),.A(I14349));
INVX1 NOT_5384 (.Y(g2608),.A(I5725));
INVX1 NOT_5385 (.Y(I9829),.A(g5013));
INVX1 NOT_5386 (.Y(I16760),.A(g10888));
INVX1 NOT_5387 (.Y(g2220),.A(g104));
INVX1 NOT_5388 (.Y(g4427),.A(g3638));
INVX1 NOT_5389 (.Y(I12930),.A(g7896));
INVX1 NOT_5390 (.Y(g7450),.A(g7148));
INVX1 NOT_5391 (.Y(I12993),.A(g8044));
INVX1 NOT_5392 (.Y(I15473),.A(g10087));
INVX1 NOT_5393 (.Y(I13290),.A(g8254));
INVX1 NOT_5394 (.Y(g2779),.A(g1974));
INVX1 NOT_5395 (.Y(I6150),.A(g2122));
INVX1 NOT_5396 (.Y(g9987),.A(I15187));
INVX1 NOT_5397 (.Y(g11541),.A(g11519));
INVX1 NOT_5398 (.Y(I17610),.A(g11549));
INVX1 NOT_5399 (.Y(I11698),.A(g7057));
INVX1 NOT_5400 (.Y(g4200),.A(I7417));
INVX1 NOT_5401 (.Y(g9771),.A(g9432));
INVX1 NOT_5402 (.Y(I12694),.A(g7374));
INVX1 NOT_5403 (.Y(I12838),.A(g7682));
INVX1 NOT_5404 (.Y(g11473),.A(I17456));
INVX1 NOT_5405 (.Y(g2023),.A(g1357));
INVX1 NOT_5406 (.Y(I10078),.A(g5729));
INVX1 NOT_5407 (.Y(I17255),.A(g11344));
INVX1 NOT_5408 (.Y(g4514),.A(g3946));
INVX1 NOT_5409 (.Y(I10598),.A(g5874));
INVX1 NOT_5410 (.Y(g5783),.A(I9377));
INVX1 NOT_5411 (.Y(g4003),.A(g3144));
INVX1 NOT_5412 (.Y(g7724),.A(I12357));
INVX1 NOT_5413 (.Y(I15359),.A(g10019));
INVX1 NOT_5414 (.Y(I6409),.A(g2356));
INVX1 NOT_5415 (.Y(g8126),.A(I12989));
INVX1 NOT_5416 (.Y(I7719),.A(g3752));
INVX1 NOT_5417 (.Y(g5112),.A(g4682));
INVX1 NOT_5418 (.Y(g7379),.A(g6863));
INVX1 NOT_5419 (.Y(g5218),.A(I8647));
INVX1 NOT_5420 (.Y(g8326),.A(I13360));
INVX1 NOT_5421 (.Y(I17188),.A(g11313));
INVX1 NOT_5422 (.Y(I17124),.A(g11232));
INVX1 NOT_5423 (.Y(g5267),.A(I8711));
INVX1 NOT_5424 (.Y(I17678),.A(g11607));
INVX1 NOT_5425 (.Y(I11427),.A(g6573));
INVX1 NOT_5426 (.Y(I12487),.A(g7723));
INVX1 NOT_5427 (.Y(I15829),.A(g10203));
INVX1 NOT_5428 (.Y(I13427),.A(g8241));
INVX1 NOT_5429 (.Y(g9892),.A(I15079));
INVX1 NOT_5430 (.Y(I8039),.A(g3506));
INVX1 NOT_5431 (.Y(I7752),.A(g3407));
INVX1 NOT_5432 (.Y(g4763),.A(g3586));
INVX1 NOT_5433 (.Y(I12502),.A(g7726));
INVX1 NOT_5434 (.Y(g4191),.A(I7390));
INVX1 NOT_5435 (.Y(I11632),.A(g6931));
INVX1 NOT_5436 (.Y(g7878),.A(g7479));
INVX1 NOT_5437 (.Y(g10850),.A(I16550));
INVX1 NOT_5438 (.Y(g8760),.A(g8670));
INVX1 NOT_5439 (.Y(g11434),.A(I17353));
INVX1 NOT_5440 (.Y(g4391),.A(g3638));
INVX1 NOT_5441 (.Y(g1989),.A(g770));
INVX1 NOT_5442 (.Y(I10322),.A(g6193));
INVX1 NOT_5443 (.Y(g7289),.A(I11543));
INVX1 NOT_5444 (.Y(g7777),.A(I12496));
INVX1 NOT_5445 (.Y(g7658),.A(I12271));
INVX1 NOT_5446 (.Y(g5401),.A(I8839));
INVX1 NOT_5447 (.Y(g3408),.A(g3108));
INVX1 NOT_5448 (.Y(I10159),.A(g5936));
INVX1 NOT_5449 (.Y(g10133),.A(g10064));
INVX1 NOT_5450 (.Y(g5676),.A(I9185));
INVX1 NOT_5451 (.Y(g2451),.A(g248));
INVX1 NOT_5452 (.Y(I10901),.A(g6620));
INVX1 NOT_5453 (.Y(g4637),.A(I8039));
INVX1 NOT_5454 (.Y(I12279),.A(g7225));
INVX1 NOT_5455 (.Y(I5348),.A(g746));
INVX1 NOT_5456 (.Y(g3336),.A(I6523));
INVX1 NOT_5457 (.Y(I15344),.A(g10025));
INVX1 NOT_5458 (.Y(g6778),.A(g5987));
INVX1 NOT_5459 (.Y(g7882),.A(g7479));
INVX1 NOT_5460 (.Y(g3768),.A(I6979));
INVX1 NOT_5461 (.Y(g10896),.A(I16650));
INVX1 NOT_5462 (.Y(I13403),.A(g8236));
INVX1 NOT_5463 (.Y(g11344),.A(I17155));
INVX1 NOT_5464 (.Y(g4307),.A(g4013));
INVX1 NOT_5465 (.Y(g4536),.A(g3880));
INVX1 NOT_5466 (.Y(g10228),.A(I15604));
INVX1 NOT_5467 (.Y(g4159),.A(I7300));
INVX1 NOT_5468 (.Y(g2346),.A(I5414));
INVX1 NOT_5469 (.Y(g4359),.A(g3880));
INVX1 NOT_5470 (.Y(I12469),.A(g7531));
INVX1 NOT_5471 (.Y(g6735),.A(I10736));
INVX1 NOT_5472 (.Y(g8183),.A(I13102));
INVX1 NOT_5473 (.Y(g8608),.A(g8482));
INVX1 NOT_5474 (.Y(g8924),.A(I14249));
INVX1 NOT_5475 (.Y(g5830),.A(I9446));
INVX1 NOT_5476 (.Y(g7611),.A(I12183));
INVX1 NOT_5477 (.Y(g8220),.A(g7826));
INVX1 NOT_5478 (.Y(I12286),.A(g7231));
INVX1 NOT_5479 (.Y(I14561),.A(g9025));
INVX1 NOT_5480 (.Y(g5727),.A(I9273));
INVX1 NOT_5481 (.Y(g2103),.A(I4961));
INVX1 NOT_5482 (.Y(I8919),.A(g4576));
INVX1 NOT_5483 (.Y(g3943),.A(g2779));
INVX1 NOT_5484 (.Y(I9177),.A(g4904));
INVX1 NOT_5485 (.Y(I7233),.A(g2817));
INVX1 NOT_5486 (.Y(I10144),.A(g5689));
INVX1 NOT_5487 (.Y(g9340),.A(I14525));
INVX1 NOT_5488 (.Y(I14295),.A(g8806));
INVX1 NOT_5489 (.Y(I9377),.A(g5576));
INVX1 NOT_5490 (.Y(I17219),.A(g11292));
INVX1 NOT_5491 (.Y(g7799),.A(I12562));
INVX1 NOT_5492 (.Y(g4757),.A(I8109));
INVX1 NOT_5493 (.Y(I16604),.A(g10786));
INVX1 NOT_5494 (.Y(I7054),.A(g3093));
INVX1 NOT_5495 (.Y(I11572),.A(g6822));
INVX1 NOT_5496 (.Y(g8423),.A(I13583));
INVX1 NOT_5497 (.Y(g6475),.A(g5987));
INVX1 NOT_5498 (.Y(g4416),.A(g3638));
INVX1 NOT_5499 (.Y(g7981),.A(g7624));
INVX1 NOT_5500 (.Y(g6949),.A(I11091));
INVX1 NOT_5501 (.Y(g3228),.A(I6409));
INVX1 NOT_5502 (.Y(g8977),.A(I14352));
INVX1 NOT_5503 (.Y(g2732),.A(I5792));
INVX1 NOT_5504 (.Y(I9287),.A(g5576));
INVX1 NOT_5505 (.Y(g9082),.A(g8892));
INVX1 NOT_5506 (.Y(g10310),.A(I15736));
INVX1 NOT_5507 (.Y(g8588),.A(I13831));
INVX1 NOT_5508 (.Y(g7997),.A(g7697));
INVX1 NOT_5509 (.Y(g2753),.A(I5827));
INVX1 NOT_5510 (.Y(I12601),.A(g7629));
INVX1 NOT_5511 (.Y(g6292),.A(I10135));
INVX1 NOT_5512 (.Y(I11127),.A(g6452));
INVX1 NOT_5513 (.Y(g4315),.A(g3863));
INVX1 NOT_5514 (.Y(g4811),.A(g3661));
INVX1 NOT_5515 (.Y(g2508),.A(g940));
INVX1 NOT_5516 (.Y(g8361),.A(I13463));
INVX1 NOT_5517 (.Y(g10379),.A(I15861));
INVX1 NOT_5518 (.Y(I10966),.A(g6561));
INVX1 NOT_5519 (.Y(g2240),.A(g88));
INVX1 NOT_5520 (.Y(I8004),.A(g3967));
INVX1 NOT_5521 (.Y(g2072),.A(I4876));
INVX1 NOT_5522 (.Y(g3433),.A(I6648));
INVX1 NOT_5523 (.Y(I6921),.A(g2839));
INVX1 NOT_5524 (.Y(I5279),.A(g73));
INVX1 NOT_5525 (.Y(g7332),.A(I11644));
INVX1 NOT_5526 (.Y(g10050),.A(I15269));
INVX1 NOT_5527 (.Y(I9199),.A(g4935));
INVX1 NOT_5528 (.Y(g10378),.A(I15858));
INVX1 NOT_5529 (.Y(I8647),.A(g4219));
INVX1 NOT_5530 (.Y(I9399),.A(g5013));
INVX1 NOT_5531 (.Y(g5624),.A(I9056));
INVX1 NOT_5532 (.Y(g7680),.A(g7148));
INVX1 NOT_5533 (.Y(g11506),.A(I17537));
INVX1 NOT_5534 (.Y(g7353),.A(I11707));
INVX1 NOT_5535 (.Y(g2043),.A(g1801));
INVX1 NOT_5536 (.Y(g6084),.A(I9731));
INVX1 NOT_5537 (.Y(g8327),.A(g8164));
INVX1 NOT_5538 (.Y(I14364),.A(g8952));
INVX1 NOT_5539 (.Y(g4874),.A(I8215));
INVX1 NOT_5540 (.Y(g6039),.A(I9652));
INVX1 NOT_5541 (.Y(g5068),.A(g4840));
INVX1 NOT_5542 (.Y(I11956),.A(g6912));
INVX1 NOT_5543 (.Y(g3096),.A(g2482));
INVX1 NOT_5544 (.Y(I13956),.A(g8451));
INVX1 NOT_5545 (.Y(I13376),.A(g8226));
INVX1 NOT_5546 (.Y(I13385),.A(g8230));
INVX1 NOT_5547 (.Y(I11103),.A(g6667));
INVX1 NOT_5548 (.Y(g3496),.A(I6686));
INVX1 NOT_5549 (.Y(g7744),.A(I12397));
INVX1 NOT_5550 (.Y(I11889),.A(g6898));
INVX1 NOT_5551 (.Y(I17470),.A(g11452));
INVX1 NOT_5552 (.Y(g7802),.A(I12571));
INVX1 NOT_5553 (.Y(I5652),.A(g554));
INVX1 NOT_5554 (.Y(g8146),.A(g8033));
INVX1 NOT_5555 (.Y(I5057),.A(g1961));
INVX1 NOT_5556 (.Y(I11354),.A(g6553));
INVX1 NOT_5557 (.Y(g2116),.A(I5020));
INVX1 NOT_5558 (.Y(g8346),.A(I13418));
INVX1 NOT_5559 (.Y(I5843),.A(g2509));
INVX1 NOT_5560 (.Y(I13354),.A(g8214));
INVX1 NOT_5561 (.Y(I8503),.A(g4445));
INVX1 NOT_5562 (.Y(I5989),.A(g2252));
INVX1 NOT_5563 (.Y(I9510),.A(g5421));
INVX1 NOT_5564 (.Y(I11824),.A(g7246));
INVX1 NOT_5565 (.Y(g2034),.A(g1766));
INVX1 NOT_5566 (.Y(g5677),.A(I9188));
INVX1 NOT_5567 (.Y(g8103),.A(g7994));
INVX1 NOT_5568 (.Y(g3395),.A(I6601));
INVX1 NOT_5569 (.Y(g2434),.A(g1362));
INVX1 NOT_5570 (.Y(g3337),.A(g2745));
INVX1 NOT_5571 (.Y(g3913),.A(g2920));
INVX1 NOT_5572 (.Y(I10289),.A(g6003));
INVX1 NOT_5573 (.Y(I17277),.A(g11390));
INVX1 NOT_5574 (.Y(I12168),.A(g7256));
INVX1 NOT_5575 (.Y(I11671),.A(g7047));
INVX1 NOT_5576 (.Y(g9310),.A(I14503));
INVX1 NOT_5577 (.Y(g6583),.A(I10535));
INVX1 NOT_5578 (.Y(g6702),.A(g5949));
INVX1 NOT_5579 (.Y(g4880),.A(g3638));
INVX1 NOT_5580 (.Y(g5866),.A(g5361));
INVX1 NOT_5581 (.Y(g8696),.A(g8656));
INVX1 NOT_5582 (.Y(I5549),.A(g868));
INVX1 NOT_5583 (.Y(I7029),.A(g2946));
INVX1 NOT_5584 (.Y(I14309),.A(g8813));
INVX1 NOT_5585 (.Y(g2347),.A(g1945));
INVX1 NOT_5586 (.Y(I7429),.A(g3344));
INVX1 NOT_5587 (.Y(g10802),.A(I16510));
INVX1 NOT_5588 (.Y(g5149),.A(I8551));
INVX1 NOT_5589 (.Y(I9144),.A(g5007));
INVX1 NOT_5590 (.Y(I14224),.A(g8794));
INVX1 NOT_5591 (.Y(g6919),.A(g6453));
INVX1 NOT_5592 (.Y(I10308),.A(g6003));
INVX1 NOT_5593 (.Y(I12363),.A(g7187));
INVX1 NOT_5594 (.Y(I7956),.A(g3428));
INVX1 NOT_5595 (.Y(g7901),.A(g7712));
INVX1 NOT_5596 (.Y(g4272),.A(g3586));
INVX1 NOT_5597 (.Y(I8320),.A(g4452));
INVX1 NOT_5598 (.Y(g10730),.A(I16407));
INVX1 NOT_5599 (.Y(I12478),.A(g7560));
INVX1 NOT_5600 (.Y(I12015),.A(g6924));
INVX1 NOT_5601 (.Y(g6276),.A(I10087));
INVX1 NOT_5602 (.Y(g11649),.A(I17749));
INVX1 NOT_5603 (.Y(g9824),.A(I14973));
INVX1 NOT_5604 (.Y(g4243),.A(g3524));
INVX1 NOT_5605 (.Y(g3266),.A(I6436));
INVX1 NOT_5606 (.Y(I9259),.A(g5301));
INVX1 NOT_5607 (.Y(g8240),.A(g7972));
INVX1 NOT_5608 (.Y(g2914),.A(I6091));
INVX1 NOT_5609 (.Y(g5198),.A(I8614));
INVX1 NOT_5610 (.Y(g5747),.A(I9317));
INVX1 NOT_5611 (.Y(I15491),.A(g10093));
INVX1 NOT_5612 (.Y(g2210),.A(g103));
INVX1 NOT_5613 (.Y(g4417),.A(I7757));
INVX1 NOT_5614 (.Y(I10495),.A(g6144));
INVX1 NOT_5615 (.Y(g8472),.A(I13666));
INVX1 NOT_5616 (.Y(g6561),.A(g5773));
INVX1 NOT_5617 (.Y(g11648),.A(I17746));
INVX1 NOT_5618 (.Y(g4935),.A(g4420));
INVX1 NOT_5619 (.Y(g9762),.A(I14903));
INVX1 NOT_5620 (.Y(I17419),.A(g11421));
INVX1 NOT_5621 (.Y(I12556),.A(g7678));
INVX1 NOT_5622 (.Y(I15604),.A(g10148));
INVX1 NOT_5623 (.Y(I10816),.A(g6406));
INVX1 NOT_5624 (.Y(I9923),.A(g5308));
INVX1 NOT_5625 (.Y(g2013),.A(g1101));
INVX1 NOT_5626 (.Y(g8443),.A(I13627));
INVX1 NOT_5627 (.Y(g7600),.A(I12150));
INVX1 NOT_5628 (.Y(I12580),.A(g7540));
INVX1 NOT_5629 (.Y(g7574),.A(g6995));
INVX1 NOT_5630 (.Y(I6085),.A(g2234));
INVX1 NOT_5631 (.Y(g10548),.A(I16209));
INVX1 NOT_5632 (.Y(I17155),.A(g11310));
INVX1 NOT_5633 (.Y(g3142),.A(I6360));
INVX1 NOT_5634 (.Y(g5241),.A(g4386));
INVX1 NOT_5635 (.Y(g6527),.A(I10445));
INVX1 NOT_5636 (.Y(I12223),.A(g7049));
INVX1 NOT_5637 (.Y(g4328),.A(g4130));
INVX1 NOT_5638 (.Y(I14687),.A(g9258));
INVX1 NOT_5639 (.Y(I17170),.A(g11294));
INVX1 NOT_5640 (.Y(I14976),.A(g9670));
INVX1 NOT_5641 (.Y(g8116),.A(I12971));
INVX1 NOT_5642 (.Y(g3255),.A(I6421));
INVX1 NOT_5643 (.Y(I7639),.A(g3722));
INVX1 NOT_5644 (.Y(g8316),.A(I13332));
INVX1 NOT_5645 (.Y(g3815),.A(g3228));
INVX1 NOT_5646 (.Y(I11211),.A(g6527));
INVX1 NOT_5647 (.Y(I10374),.A(g5852));
INVX1 NOT_5648 (.Y(g6764),.A(g5987));
INVX1 NOT_5649 (.Y(I7109),.A(g2970));
INVX1 NOT_5650 (.Y(I5909),.A(g2207));
INVX1 NOT_5651 (.Y(I16534),.A(g10747));
INVX1 NOT_5652 (.Y(I10643),.A(g6026));
INVX1 NOT_5653 (.Y(I11088),.A(g6434));
INVX1 NOT_5654 (.Y(I11024),.A(g6399));
INVX1 NOT_5655 (.Y(g9556),.A(I14701));
INVX1 NOT_5656 (.Y(I16098),.A(g10369));
INVX1 NOT_5657 (.Y(g10317),.A(I15749));
INVX1 NOT_5658 (.Y(g8565),.A(I13788));
INVX1 NOT_5659 (.Y(g2820),.A(I5926));
INVX1 NOT_5660 (.Y(g3097),.A(g2482));
INVX1 NOT_5661 (.Y(I9886),.A(g5286));
INVX1 NOT_5662 (.Y(I6941),.A(g2858));
INVX1 NOT_5663 (.Y(g3726),.A(I6898));
INVX1 NOT_5664 (.Y(g7580),.A(I12056));
INVX1 NOT_5665 (.Y(g6503),.A(I10421));
INVX1 NOT_5666 (.Y(g5644),.A(I9093));
INVX1 NOT_5667 (.Y(I5740),.A(g2341));
INVX1 NOT_5668 (.Y(g6970),.A(I11122));
INVX1 NOT_5669 (.Y(g8347),.A(I13421));
INVX1 NOT_5670 (.Y(I15395),.A(g10058));
INVX1 NOT_5671 (.Y(g2317),.A(g622));
INVX1 NOT_5672 (.Y(I8892),.A(g4554));
INVX1 NOT_5673 (.Y(g10129),.A(I15389));
INVX1 NOT_5674 (.Y(g9930),.A(I15127));
INVX1 NOT_5675 (.Y(I9114),.A(g5603));
INVX1 NOT_5676 (.Y(g6925),.A(I11043));
INVX1 NOT_5677 (.Y(I17194),.A(g11317));
INVX1 NOT_5678 (.Y(I7707),.A(g3370));
INVX1 NOT_5679 (.Y(g11395),.A(I17228));
INVX1 NOT_5680 (.Y(g1962),.A(g27));
INVX1 NOT_5681 (.Y(g10057),.A(I15278));
INVX1 NOT_5682 (.Y(g2601),.A(I5704));
INVX1 NOT_5683 (.Y(g10128),.A(I15386));
INVX1 NOT_5684 (.Y(g5818),.A(g5320));
INVX1 NOT_5685 (.Y(g8697),.A(g8660));
INVX1 NOT_5686 (.Y(I6520),.A(g3186));
INVX1 NOT_5687 (.Y(I14668),.A(g9309));
INVX1 NOT_5688 (.Y(g4213),.A(I7456));
INVX1 NOT_5689 (.Y(g11633),.A(I17713));
INVX1 NOT_5690 (.Y(I11659),.A(g7097));
INVX1 NOT_5691 (.Y(I12186),.A(g7264));
INVX1 NOT_5692 (.Y(g6120),.A(I9813));
INVX1 NOT_5693 (.Y(I10195),.A(g6116));
INVX1 NOT_5694 (.Y(I6031),.A(g2209));
INVX1 NOT_5695 (.Y(I12953),.A(g8024));
INVX1 NOT_5696 (.Y(g10323),.A(I15763));
INVX1 NOT_5697 (.Y(g11191),.A(g11112));
INVX1 NOT_5698 (.Y(g2775),.A(I5862));
INVX1 NOT_5699 (.Y(g7076),.A(I11303));
INVX1 NOT_5700 (.Y(I6812),.A(g3290));
INVX1 NOT_5701 (.Y(g3783),.A(I7009));
INVX1 NOT_5702 (.Y(g7476),.A(g6933));
INVX1 NOT_5703 (.Y(I6958),.A(g2872));
INVX1 NOT_5704 (.Y(g5893),.A(g5106));
INVX1 NOT_5705 (.Y(g6277),.A(I10090));
INVX1 NOT_5706 (.Y(I14525),.A(g9109));
INVX1 NOT_5707 (.Y(I14424),.A(g8945));
INVX1 NOT_5708 (.Y(g3112),.A(g2482));
INVX1 NOT_5709 (.Y(g3267),.A(I6439));
INVX1 NOT_5710 (.Y(g10775),.A(I16461));
INVX1 NOT_5711 (.Y(I16766),.A(g10892));
INVX1 NOT_5712 (.Y(I12936),.A(g7983));
INVX1 NOT_5713 (.Y(I15832),.A(g10206));
INVX1 NOT_5714 (.Y(I8340),.A(g4804));
INVX1 NOT_5715 (.Y(I11296),.A(g6525));
INVX1 NOT_5716 (.Y(g2060),.A(g1380));
INVX1 NOT_5717 (.Y(g6617),.A(g6019));
INVX1 NOT_5718 (.Y(I14558),.A(g9024));
INVX1 NOT_5719 (.Y(g6789),.A(I10789));
INVX1 NOT_5720 (.Y(I17749),.A(g11644));
INVX1 NOT_5721 (.Y(I11644),.A(g6970));
INVX1 NOT_5722 (.Y(I17616),.A(g11561));
INVX1 NOT_5723 (.Y(I16871),.A(g10973));
INVX1 NOT_5724 (.Y(I11338),.A(g6680));
INVX1 NOT_5725 (.Y(I13338),.A(g8210));
INVX1 NOT_5726 (.Y(I9594),.A(g5083));
INVX1 NOT_5727 (.Y(g4166),.A(I7315));
INVX1 NOT_5728 (.Y(g11440),.A(I17371));
INVX1 NOT_5729 (.Y(g4366),.A(I7659));
INVX1 NOT_5730 (.Y(g5426),.A(I8869));
INVX1 NOT_5731 (.Y(I15861),.A(g10339));
INVX1 NOT_5732 (.Y(I16360),.A(g10590));
INVX1 NOT_5733 (.Y(I6911),.A(g2825));
INVX1 NOT_5734 (.Y(I13969),.A(g8451));
INVX1 NOT_5735 (.Y(I7833),.A(g3585));
INVX1 NOT_5736 (.Y(g7285),.A(I11531));
INVX1 NOT_5737 (.Y(g3329),.A(I6504));
INVX1 NOT_5738 (.Y(I15247),.A(g10032));
INVX1 NOT_5739 (.Y(g11573),.A(g11561));
INVX1 NOT_5740 (.Y(I5525),.A(g589));
INVX1 NOT_5741 (.Y(I5710),.A(g2431));
INVX1 NOT_5742 (.Y(g3761),.A(I6962));
INVX1 NOT_5743 (.Y(g5614),.A(I9040));
INVX1 NOT_5744 (.Y(I12762),.A(g7541));
INVX1 NOT_5745 (.Y(I17704),.A(g11618));
INVX1 NOT_5746 (.Y(g4056),.A(I7173));
INVX1 NOT_5747 (.Y(g7500),.A(g6943));
INVX1 NOT_5748 (.Y(I10713),.A(g6003));
INVX1 NOT_5749 (.Y(g8317),.A(I13335));
INVX1 NOT_5750 (.Y(I15389),.A(g10110));
INVX1 NOT_5751 (.Y(g4456),.A(g3375));
INVX1 NOT_5752 (.Y(I14713),.A(g9052));
INVX1 NOT_5753 (.Y(g6299),.A(I10156));
INVX1 NOT_5754 (.Y(g5821),.A(I9433));
INVX1 NOT_5755 (.Y(g3828),.A(g2920));
INVX1 NOT_5756 (.Y(g10697),.A(I16370));
INVX1 NOT_5757 (.Y(g6547),.A(g5893));
INVX1 NOT_5758 (.Y(I13197),.A(g8186));
INVX1 NOT_5759 (.Y(g11389),.A(I17216));
INVX1 NOT_5760 (.Y(g11045),.A(I16796));
INVX1 NOT_5761 (.Y(I6733),.A(g3321));
INVX1 NOT_5762 (.Y(I9065),.A(g4760));
INVX1 NOT_5763 (.Y(I17466),.A(g11447));
INVX1 NOT_5764 (.Y(g8601),.A(g8477));
INVX1 NOT_5765 (.Y(g10261),.A(g10126));
INVX1 NOT_5766 (.Y(g2937),.A(I6106));
INVX1 NOT_5767 (.Y(g3727),.A(I6901));
INVX1 NOT_5768 (.Y(g2079),.A(I4891));
INVX1 NOT_5769 (.Y(g5984),.A(I9602));
INVX1 NOT_5770 (.Y(I10610),.A(g5879));
INVX1 NOT_5771 (.Y(g10880),.A(I16610));
INVX1 NOT_5772 (.Y(I15701),.A(g10236));
INVX1 NOT_5773 (.Y(g4355),.A(I7642));
INVX1 NOT_5774 (.Y(g11388),.A(I17213));
INVX1 NOT_5775 (.Y(g7339),.A(I11665));
INVX1 NOT_5776 (.Y(g2479),.A(g26));
INVX1 NOT_5777 (.Y(I10042),.A(g5723));
INVX1 NOT_5778 (.Y(I15272),.A(g10019));
INVX1 NOT_5779 (.Y(I16629),.A(g10860));
INVX1 NOT_5780 (.Y(g2840),.A(I5960));
INVX1 NOT_5781 (.Y(I10189),.A(g6112));
INVX1 NOT_5782 (.Y(g7024),.A(I11169));
INVX1 NOT_5783 (.Y(I16220),.A(g10502));
INVX1 NOT_5784 (.Y(g2190),.A(I5149));
INVX1 NOT_5785 (.Y(g4260),.A(I7513));
INVX1 NOT_5786 (.Y(g2390),.A(I5475));
INVX1 NOT_5787 (.Y(g7795),.A(I12550));
INVX1 NOT_5788 (.Y(I9433),.A(g5069));
INVX1 NOT_5789 (.Y(I17642),.A(g11579));
INVX1 NOT_5790 (.Y(I10678),.A(g5777));
INVX1 NOT_5791 (.Y(g7737),.A(I12388));
INVX1 NOT_5792 (.Y(g7809),.A(I12592));
INVX1 NOT_5793 (.Y(g3703),.A(g2920));
INVX1 NOT_5794 (.Y(I14188),.A(g8792));
INVX1 NOT_5795 (.Y(I14678),.A(g9265));
INVX1 NOT_5796 (.Y(g5106),.A(I8490));
INVX1 NOT_5797 (.Y(g4463),.A(g3829));
INVX1 NOT_5798 (.Y(I9096),.A(g5568));
INVX1 NOT_5799 (.Y(g2156),.A(I5073));
INVX1 NOT_5800 (.Y(g7672),.A(I12293));
INVX1 NOT_5801 (.Y(I14939),.A(g9454));
INVX1 NOT_5802 (.Y(g2356),.A(I5438));
INVX1 NOT_5803 (.Y(g7077),.A(I11306));
INVX1 NOT_5804 (.Y(g6709),.A(g5949));
INVX1 NOT_5805 (.Y(I17733),.A(g11639));
INVX1 NOT_5806 (.Y(g9814),.A(g9490));
INVX1 NOT_5807 (.Y(g5790),.A(I9388));
INVX1 NOT_5808 (.Y(I9550),.A(g5030));
INVX1 NOT_5809 (.Y(I10030),.A(g5685));
INVX1 NOT_5810 (.Y(g7477),.A(I11869));
INVX1 NOT_5811 (.Y(I10093),.A(g5779));
INVX1 NOT_5812 (.Y(I9845),.A(g5405));
INVX1 NOT_5813 (.Y(g3624),.A(I6767));
INVX1 NOT_5814 (.Y(g6140),.A(I9851));
INVX1 NOT_5815 (.Y(g6340),.A(I10243));
INVX1 NOT_5816 (.Y(I5111),.A(g39));
INVX1 NOT_5817 (.Y(I11581),.A(g6826));
INVX1 NOT_5818 (.Y(I11450),.A(g6488));
INVX1 NOT_5819 (.Y(I12568),.A(g7502));
INVX1 NOT_5820 (.Y(g9350),.A(I14555));
INVX1 NOT_5821 (.Y(g10499),.A(I16124));
INVX1 NOT_5822 (.Y(I5311),.A(g98));
INVX1 NOT_5823 (.Y(g3068),.A(g2303));
INVX1 NOT_5824 (.Y(I13714),.A(g8351));
INVX1 NOT_5825 (.Y(I11315),.A(g6644));
INVX1 NOT_5826 (.Y(g8784),.A(I14087));
INVX1 NOT_5827 (.Y(g2942),.A(I6121));
INVX1 NOT_5828 (.Y(g8739),.A(g8640));
INVX1 NOT_5829 (.Y(I12242),.A(g7089));
INVX1 NOT_5830 (.Y(g4279),.A(I7536));
INVX1 NOT_5831 (.Y(I11707),.A(g7009));
INVX1 NOT_5832 (.Y(g7205),.A(I11433));
INVX1 NOT_5833 (.Y(g9773),.A(g9474));
INVX1 NOT_5834 (.Y(I7086),.A(g3142));
INVX1 NOT_5835 (.Y(I13819),.A(g8488));
INVX1 NOT_5836 (.Y(g11061),.A(g10974));
INVX1 NOT_5837 (.Y(g10498),.A(I16121));
INVX1 NOT_5838 (.Y(g9009),.A(I14405));
INVX1 NOT_5839 (.Y(g6435),.A(I10355));
INVX1 NOT_5840 (.Y(g4167),.A(I7318));
INVX1 NOT_5841 (.Y(g5027),.A(I8396));
INVX1 NOT_5842 (.Y(g6517),.A(I10434));
INVX1 NOT_5843 (.Y(g6082),.A(I9727));
INVX1 NOT_5844 (.Y(I12123),.A(g6861));
INVX1 NOT_5845 (.Y(g4318),.A(g4130));
INVX1 NOT_5846 (.Y(g4367),.A(I7662));
INVX1 NOT_5847 (.Y(I16859),.A(g10911));
INVX1 NOT_5848 (.Y(g4872),.A(I8211));
INVX1 NOT_5849 (.Y(g7634),.A(I12242));
INVX1 NOT_5850 (.Y(I5174),.A(g52));
INVX1 NOT_5851 (.Y(I16950),.A(g11081));
INVX1 NOT_5852 (.Y(g8079),.A(I12939));
INVX1 NOT_5853 (.Y(I16370),.A(g10592));
INVX1 NOT_5854 (.Y(g6482),.A(I10412));
INVX1 NOT_5855 (.Y(I11055),.A(g6419));
INVX1 NOT_5856 (.Y(g10056),.A(I15275));
INVX1 NOT_5857 (.Y(I9807),.A(g5419));
INVX1 NOT_5858 (.Y(g8479),.A(g8319));
INVX1 NOT_5859 (.Y(I7185),.A(g2626));
INVX1 NOT_5860 (.Y(I12751),.A(g7626));
INVX1 NOT_5861 (.Y(g9769),.A(I14918));
INVX1 NOT_5862 (.Y(g4057),.A(I7176));
INVX1 NOT_5863 (.Y(g5904),.A(I9539));
INVX1 NOT_5864 (.Y(g7304),.A(I11560));
INVX1 NOT_5865 (.Y(g5200),.A(g4567));
INVX1 NOT_5866 (.Y(g10080),.A(I15308));
INVX1 NOT_5867 (.Y(g8294),.A(I13236));
INVX1 NOT_5868 (.Y(I13978),.A(g8575));
INVX1 NOT_5869 (.Y(g4457),.A(g3829));
INVX1 NOT_5870 (.Y(g2163),.A(I5092));
INVX1 NOT_5871 (.Y(I8877),.A(g4421));
INVX1 NOT_5872 (.Y(g2363),.A(I5441));
INVX1 NOT_5873 (.Y(I7070),.A(g3138));
INVX1 NOT_5874 (.Y(g5446),.A(I8877));
INVX1 NOT_5875 (.Y(I11590),.A(g6829));
INVX1 NOT_5876 (.Y(I16172),.A(g10498));
INVX1 NOT_5877 (.Y(g4193),.A(I7396));
INVX1 NOT_5878 (.Y(g3716),.A(I6876));
INVX1 NOT_5879 (.Y(g11360),.A(I17185));
INVX1 NOT_5880 (.Y(g4393),.A(I7726));
INVX1 NOT_5881 (.Y(I10837),.A(g6717));
INVX1 NOT_5882 (.Y(g2432),.A(I5513));
INVX1 NOT_5883 (.Y(I12293),.A(g7116));
INVX1 NOT_5884 (.Y(g10271),.A(I15665));
INVX1 NOT_5885 (.Y(I12638),.A(g7708));
INVX1 NOT_5886 (.Y(g11447),.A(I17390));
INVX1 NOT_5887 (.Y(I13741),.A(g8296));
INVX1 NOT_5888 (.Y(I15162),.A(g9958));
INVX1 NOT_5889 (.Y(g4549),.A(I7956));
INVX1 NOT_5890 (.Y(I17555),.A(g11503));
INVX1 NOT_5891 (.Y(I6898),.A(g2964));
INVX1 NOT_5892 (.Y(I12265),.A(g7211));
INVX1 NOT_5893 (.Y(g11162),.A(g10950));
INVX1 NOT_5894 (.Y(g7754),.A(I12427));
INVX1 NOT_5895 (.Y(g10461),.A(I15974));
INVX1 NOT_5896 (.Y(g5191),.A(g4640));
INVX1 NOT_5897 (.Y(g8156),.A(I13051));
INVX1 NOT_5898 (.Y(I9248),.A(g4954));
INVX1 NOT_5899 (.Y(g3747),.A(g3015));
INVX1 NOT_5900 (.Y(I11094),.A(g6657));
INVX1 NOT_5901 (.Y(g1973),.A(g466));
INVX1 NOT_5902 (.Y(g5391),.A(I8827));
INVX1 NOT_5903 (.Y(g8356),.A(I13448));
INVX1 NOT_5904 (.Y(g10342),.A(I15792));
INVX1 NOT_5905 (.Y(g3398),.A(g2896));
INVX1 NOT_5906 (.Y(g6214),.A(g5446));
INVX1 NOT_5907 (.Y(g7273),.A(g6365));
INVX1 NOT_5908 (.Y(I5020),.A(g1176));
INVX1 NOT_5909 (.Y(I6510),.A(g3267));
INVX1 NOT_5910 (.Y(g9993),.A(I15193));
INVX1 NOT_5911 (.Y(g10145),.A(I15437));
INVX1 NOT_5912 (.Y(g10031),.A(I15229));
INVX1 NOT_5913 (.Y(g6110),.A(I9783));
INVX1 NOT_5914 (.Y(g5637),.A(I9074));
INVX1 NOT_5915 (.Y(g6310),.A(I10189));
INVX1 NOT_5916 (.Y(g11629),.A(I17701));
INVX1 NOT_5917 (.Y(g9822),.A(I14967));
INVX1 NOT_5918 (.Y(g10199),.A(g10172));
INVX1 NOT_5919 (.Y(g11451),.A(I17410));
INVX1 NOT_5920 (.Y(g11472),.A(I17453));
INVX1 NOT_5921 (.Y(g7044),.A(I11217));
INVX1 NOT_5922 (.Y(g10887),.A(I16623));
INVX1 NOT_5923 (.Y(g2912),.A(I6085));
INVX1 NOT_5924 (.Y(I13735),.A(g8293));
INVX1 NOT_5925 (.Y(g1969),.A(g456));
INVX1 NOT_5926 (.Y(g4121),.A(I7264));
INVX1 NOT_5927 (.Y(g5107),.A(g4459));
INVX1 NOT_5928 (.Y(g8704),.A(g8667));
INVX1 NOT_5929 (.Y(g4321),.A(g3863));
INVX1 NOT_5930 (.Y(g2157),.A(g1703));
INVX1 NOT_5931 (.Y(g11628),.A(I17698));
INVX1 NOT_5932 (.Y(g10198),.A(I15568));
INVX1 NOT_5933 (.Y(I7131),.A(g2640));
INVX1 NOT_5934 (.Y(I7006),.A(g2912));
INVX1 NOT_5935 (.Y(g7983),.A(I12793));
INVX1 NOT_5936 (.Y(I10201),.A(g5998));
INVX1 NOT_5937 (.Y(g5223),.A(g4640));
INVX1 NOT_5938 (.Y(I11695),.A(g7052));
INVX1 NOT_5939 (.Y(g10528),.A(g10464));
INVX1 NOT_5940 (.Y(g10696),.A(g10621));
INVX1 NOT_5941 (.Y(g4232),.A(I7487));
INVX1 NOT_5942 (.Y(I12835),.A(g7660));
INVX1 NOT_5943 (.Y(I13695),.A(g8363));
INVX1 NOT_5944 (.Y(g10330),.A(I15778));
INVX1 NOT_5945 (.Y(g5858),.A(I9475));
INVX1 NOT_5946 (.Y(g10393),.A(g10317));
INVX1 NOT_5947 (.Y(I10075),.A(g5724));
INVX1 NOT_5948 (.Y(I7766),.A(g3770));
INVX1 NOT_5949 (.Y(g8954),.A(I14315));
INVX1 NOT_5950 (.Y(I16540),.A(g10722));
INVX1 NOT_5951 (.Y(g6236),.A(I9981));
INVX1 NOT_5952 (.Y(I6694),.A(g2749));
INVX1 NOT_5953 (.Y(g7543),.A(I11961));
INVX1 NOT_5954 (.Y(I12586),.A(g7561));
INVX1 NOT_5955 (.Y(g11071),.A(g10913));
INVX1 NOT_5956 (.Y(g8363),.A(I13469));
INVX1 NOT_5957 (.Y(I7487),.A(g3371));
INVX1 NOT_5958 (.Y(I8237),.A(g4295));
INVX1 NOT_5959 (.Y(g5416),.A(I8851));
INVX1 NOT_5960 (.Y(I14494),.A(g8887));
INVX1 NOT_5961 (.Y(g3119),.A(I6347));
INVX1 NOT_5962 (.Y(g10132),.A(g10063));
INVX1 NOT_5963 (.Y(I17519),.A(g11484));
INVX1 NOT_5964 (.Y(g10869),.A(I16577));
INVX1 NOT_5965 (.Y(I6088),.A(g2235));
INVX1 NOT_5966 (.Y(I17176),.A(g11286));
INVX1 NOT_5967 (.Y(I17185),.A(g11311));
INVX1 NOT_5968 (.Y(I10623),.A(g6002));
INVX1 NOT_5969 (.Y(I12442),.A(g7672));
INVX1 NOT_5970 (.Y(I17675),.A(g11606));
INVX1 NOT_5971 (.Y(I17092),.A(g11217));
INVX1 NOT_5972 (.Y(I16203),.A(g10454));
INVX1 NOT_5973 (.Y(g4519),.A(I7920));
INVX1 NOT_5974 (.Y(g5251),.A(g4640));
INVX1 NOT_5975 (.Y(g6590),.A(g5949));
INVX1 NOT_5976 (.Y(g6877),.A(I10963));
INVX1 NOT_5977 (.Y(I4777),.A(g18));
INVX1 NOT_5978 (.Y(g10868),.A(I16574));
INVX1 NOT_5979 (.Y(g5811),.A(I9415));
INVX1 NOT_5980 (.Y(g5642),.A(I9087));
INVX1 NOT_5981 (.Y(g3352),.A(I6538));
INVX1 NOT_5982 (.Y(I9783),.A(g5395));
INVX1 NOT_5983 (.Y(g2626),.A(g2000));
INVX1 NOT_5984 (.Y(g7534),.A(I11942));
INVX1 NOT_5985 (.Y(g7729),.A(I12372));
INVX1 NOT_5986 (.Y(g7961),.A(g7664));
INVX1 NOT_5987 (.Y(g5047),.A(g4354));
INVX1 NOT_5988 (.Y(I13457),.A(g8184));
INVX1 NOT_5989 (.Y(I10984),.A(g6757));
INVX1 NOT_5990 (.Y(g9895),.A(I15088));
INVX1 NOT_5991 (.Y(g6657),.A(I10620));
INVX1 NOT_5992 (.Y(g10161),.A(I15479));
INVX1 NOT_5993 (.Y(g4552),.A(g3880));
INVX1 NOT_5994 (.Y(g4606),.A(g3829));
INVX1 NOT_5995 (.Y(I15858),.A(g10336));
INVX1 NOT_5996 (.Y(g8568),.A(I13797));
INVX1 NOT_5997 (.Y(I8089),.A(g3545));
INVX1 NOT_5998 (.Y(I10352),.A(g6216));
INVX1 NOT_5999 (.Y(g6556),.A(g5747));
INVX1 NOT_6000 (.Y(I14352),.A(g8946));
INVX1 NOT_6001 (.Y(g7927),.A(g7500));
INVX1 NOT_6002 (.Y(I10822),.A(g6584));
INVX1 NOT_6003 (.Y(g5874),.A(I9491));
INVX1 NOT_6004 (.Y(I9001),.A(g4762));
INVX1 NOT_6005 (.Y(g10259),.A(g10141));
INVX1 NOT_6006 (.Y(I14418),.A(g8941));
INVX1 NOT_6007 (.Y(g10708),.A(I16387));
INVX1 NOT_6008 (.Y(I16739),.A(g10856));
INVX1 NOT_6009 (.Y(I12430),.A(g7649));
INVX1 NOT_6010 (.Y(g3186),.A(I6373));
INVX1 NOT_6011 (.Y(g5654),.A(I9123));
INVX1 NOT_6012 (.Y(I12493),.A(g7650));
INVX1 NOT_6013 (.Y(g10471),.A(g10378));
INVX1 NOT_6014 (.Y(g7414),.A(I11794));
INVX1 NOT_6015 (.Y(I9293),.A(g5486));
INVX1 NOT_6016 (.Y(g3386),.A(g3144));
INVX1 NOT_6017 (.Y(g10087),.A(I15314));
INVX1 NOT_6018 (.Y(g8357),.A(I13451));
INVX1 NOT_6019 (.Y(I9129),.A(g4892));
INVX1 NOT_6020 (.Y(g7946),.A(g7416));
INVX1 NOT_6021 (.Y(g10258),.A(g10198));
INVX1 NOT_6022 (.Y(g3975),.A(g3121));
INVX1 NOT_6023 (.Y(I7173),.A(g2644));
INVX1 NOT_6024 (.Y(I9329),.A(g5504));
INVX1 NOT_6025 (.Y(I5973),.A(g2247));
INVX1 NOT_6026 (.Y(g4586),.A(g4089));
INVX1 NOT_6027 (.Y(g11394),.A(I17225));
INVX1 NOT_6028 (.Y(g6464),.A(I10398));
INVX1 NOT_6029 (.Y(g7903),.A(g7446));
INVX1 NOT_6030 (.Y(g2683),.A(g2037));
INVX1 NOT_6031 (.Y(I11689),.A(g7044));
INVX1 NOT_6032 (.Y(I6870),.A(g2852));
INVX1 NOT_6033 (.Y(g3274),.A(I6454));
INVX1 NOT_6034 (.Y(g3426),.A(g3121));
INVX1 NOT_6035 (.Y(g5880),.A(g5361));
INVX1 NOT_6036 (.Y(I12035),.A(g6930));
INVX1 NOT_6037 (.Y(I13280),.A(g8250));
INVX1 NOT_6038 (.Y(g2778),.A(g2276));
INVX1 NOT_6039 (.Y(g10244),.A(g10131));
INVX1 NOT_6040 (.Y(I9727),.A(g5250));
INVX1 NOT_6041 (.Y(I7369),.A(g4051));
INVX1 NOT_6042 (.Y(g3370),.A(I6560));
INVX1 NOT_6043 (.Y(I10589),.A(g5763));
INVX1 NOT_6044 (.Y(I13624),.A(g8320));
INVX1 NOT_6045 (.Y(I14194),.A(g8798));
INVX1 NOT_6046 (.Y(g11420),.A(I17315));
INVX1 NOT_6047 (.Y(g6563),.A(g5783));
INVX1 NOT_6048 (.Y(I7920),.A(g3440));
INVX1 NOT_6049 (.Y(g5272),.A(I8724));
INVX1 NOT_6050 (.Y(g11319),.A(I17116));
INVX1 NOT_6051 (.Y(g7036),.A(g6420));
INVX1 NOT_6052 (.Y(g9085),.A(g8892));
INVX1 NOT_6053 (.Y(g10069),.A(I15296));
INVX1 NOT_6054 (.Y(I7459),.A(g3720));
INVX1 NOT_6055 (.Y(I9221),.A(g5236));
INVX1 NOT_6056 (.Y(g4525),.A(g3880));
INVX1 NOT_6057 (.Y(g7436),.A(g7227));
INVX1 NOT_6058 (.Y(g8626),.A(g8498));
INVX1 NOT_6059 (.Y(g6295),.A(I10144));
INVX1 NOT_6060 (.Y(I12517),.A(g7737));
INVX1 NOT_6061 (.Y(I13102),.A(g7928));
INVX1 NOT_6062 (.Y(g6237),.A(I9984));
INVX1 NOT_6063 (.Y(g11446),.A(I17387));
INVX1 NOT_6064 (.Y(g10774),.A(I16458));
INVX1 NOT_6065 (.Y(I17438),.A(g11444));
INVX1 NOT_6066 (.Y(I10477),.A(g6049));
INVX1 NOT_6067 (.Y(I16366),.A(g10591));
INVX1 NOT_6068 (.Y(g5417),.A(I8854));
INVX1 NOT_6069 (.Y(g2075),.A(I4883));
INVX1 NOT_6070 (.Y(I14477),.A(g8943));
INVX1 NOT_6071 (.Y(g10879),.A(I16607));
INVX1 NOT_6072 (.Y(I16632),.A(g10861));
INVX1 NOT_6073 (.Y(g11059),.A(g10974));
INVX1 NOT_6074 (.Y(g6844),.A(I10904));
INVX1 NOT_6075 (.Y(g7335),.A(I11653));
INVX1 NOT_6076 (.Y(g2475),.A(g192));
INVX1 NOT_6077 (.Y(I14119),.A(g8779));
INVX1 NOT_6078 (.Y(g1988),.A(g766));
INVX1 NOT_6079 (.Y(g3544),.A(g3164));
INVX1 NOT_6080 (.Y(g2949),.A(I6150));
INVX1 NOT_6081 (.Y(g7288),.A(I11540));
INVX1 NOT_6082 (.Y(g11540),.A(g11519));
INVX1 NOT_6083 (.Y(g5982),.A(I9598));
INVX1 NOT_6084 (.Y(g10878),.A(I16604));
INVX1 NOT_6085 (.Y(I7793),.A(g3783));
INVX1 NOT_6086 (.Y(I10864),.A(g6634));
INVX1 NOT_6087 (.Y(g3636),.A(I6815));
INVX1 NOT_6088 (.Y(g5629),.A(I9065));
INVX1 NOT_6089 (.Y(I9953),.A(g5484));
INVX1 NOT_6090 (.Y(g6089),.A(g4977));
INVX1 NOT_6091 (.Y(I12193),.A(g7270));
INVX1 NOT_6092 (.Y(g10171),.A(I15507));
INVX1 NOT_6093 (.Y(g6731),.A(g6001));
INVX1 NOT_6094 (.Y(I9068),.A(g4768));
INVX1 NOT_6095 (.Y(g7805),.A(I12580));
INVX1 NOT_6096 (.Y(I5655),.A(g557));
INVX1 NOT_6097 (.Y(g7916),.A(g7651));
INVX1 NOT_6098 (.Y(g11203),.A(g11112));
INVX1 NOT_6099 (.Y(g5542),.A(I8967));
INVX1 NOT_6100 (.Y(g7022),.A(g6389));
INVX1 NOT_6101 (.Y(g3306),.A(I6477));
INVX1 NOT_6102 (.Y(g2998),.A(g2462));
INVX1 NOT_6103 (.Y(g2646),.A(g1992));
INVX1 NOT_6104 (.Y(g4158),.A(g3304));
INVX1 NOT_6105 (.Y(g7422),.A(I11810));
INVX1 NOT_6106 (.Y(g7749),.A(I12412));
INVX1 NOT_6107 (.Y(I6065),.A(g2226));
INVX1 NOT_6108 (.Y(g6557),.A(g5748));
INVX1 NOT_6109 (.Y(I12165),.A(g6882));
INVX1 NOT_6110 (.Y(I12523),.A(g7421));
INVX1 NOT_6111 (.Y(g10792),.A(I16492));
INVX1 NOT_6112 (.Y(g11044),.A(I16793));
INVX1 NOT_6113 (.Y(g3790),.A(g3228));
INVX1 NOT_6114 (.Y(I15281),.A(g10025));
INVX1 NOT_6115 (.Y(g2084),.A(I4900));
INVX1 NOT_6116 (.Y(g2603),.A(I5710));
INVX1 NOT_6117 (.Y(I8967),.A(g4482));
INVX1 NOT_6118 (.Y(g6705),.A(I10682));
INVX1 NOT_6119 (.Y(g2039),.A(g1781));
INVX1 NOT_6120 (.Y(I9677),.A(g5190));
INVX1 NOT_6121 (.Y(g3387),.A(I6587));
INVX1 NOT_6122 (.Y(I10305),.A(g6180));
INVX1 NOT_6123 (.Y(g5800),.A(I9402));
INVX1 NOT_6124 (.Y(I5410),.A(g901));
INVX1 NOT_6125 (.Y(g3461),.A(I6671));
INVX1 NOT_6126 (.Y(I15377),.A(g10104));
INVX1 NOT_6127 (.Y(g6242),.A(I9995));
INVX1 NOT_6128 (.Y(g2850),.A(I5976));
INVX1 NOT_6129 (.Y(g9431),.A(g9085));
INVX1 NOT_6130 (.Y(g7798),.A(I12559));
INVX1 NOT_6131 (.Y(g11301),.A(I17084));
INVX1 NOT_6132 (.Y(g10459),.A(I15968));
INVX1 NOT_6133 (.Y(g9812),.A(g9490));
INVX1 NOT_6134 (.Y(g3756),.A(g3015));
INVX1 NOT_6135 (.Y(g4587),.A(g3829));
INVX1 NOT_6136 (.Y(I12475),.A(g7545));
INVX1 NOT_6137 (.Y(g11377),.A(I17202));
INVX1 NOT_6138 (.Y(I9866),.A(g5274));
INVX1 NOT_6139 (.Y(g6948),.A(I11088));
INVX1 NOT_6140 (.Y(g3622),.A(I6757));
INVX1 NOT_6141 (.Y(g9958),.A(I15157));
INVX1 NOT_6142 (.Y(g7560),.A(I12012));
INVX1 NOT_6143 (.Y(g4275),.A(g3664));
INVX1 NOT_6144 (.Y(g4311),.A(g4130));
INVX1 NOT_6145 (.Y(g10458),.A(I15965));
INVX1 NOT_6146 (.Y(g8782),.A(I14083));
INVX1 NOT_6147 (.Y(g3427),.A(g3144));
INVX1 NOT_6148 (.Y(I15562),.A(g10098));
INVX1 NOT_6149 (.Y(I9349),.A(g5515));
INVX1 NOT_6150 (.Y(g6955),.A(I11103));
INVX1 NOT_6151 (.Y(I10036),.A(g5701));
INVX1 NOT_6152 (.Y(g4615),.A(I8024));
INVX1 NOT_6153 (.Y(g5213),.A(g4640));
INVX1 NOT_6154 (.Y(g11645),.A(I17739));
INVX1 NOT_6155 (.Y(I10177),.A(g6103));
INVX1 NOT_6156 (.Y(I10560),.A(g5887));
INVX1 NOT_6157 (.Y(I11456),.A(g6440));
INVX1 NOT_6158 (.Y(I14101),.A(g8774));
INVX1 NOT_6159 (.Y(I9848),.A(g5557));
INVX1 NOT_6160 (.Y(I15290),.A(g9984));
INVX1 NOT_6161 (.Y(g6254),.A(I10021));
INVX1 NOT_6162 (.Y(g8475),.A(g8314));
INVX1 NOT_6163 (.Y(g4174),.A(I7339));
INVX1 NOT_6164 (.Y(g6814),.A(I10852));
INVX1 NOT_6165 (.Y(g9765),.A(I14910));
INVX1 NOT_6166 (.Y(I17636),.A(g11577));
INVX1 NOT_6167 (.Y(I15698),.A(g10235));
INVX1 NOT_6168 (.Y(g10545),.A(I16200));
INVX1 NOT_6169 (.Y(g2919),.A(I6102));
INVX1 NOT_6170 (.Y(g7037),.A(I11198));
INVX1 NOT_6171 (.Y(g10079),.A(I15305));
INVX1 NOT_6172 (.Y(g10444),.A(g10325));
INVX1 NOT_6173 (.Y(I9699),.A(g5426));
INVX1 NOT_6174 (.Y(g6150),.A(I9869));
INVX1 NOT_6175 (.Y(I14642),.A(g9088));
INVX1 NOT_6176 (.Y(g7437),.A(I11829));
INVX1 NOT_6177 (.Y(I16784),.A(g10895));
INVX1 NOT_6178 (.Y(I5667),.A(g566));
INVX1 NOT_6179 (.Y(I6395),.A(g2334));
INVX1 NOT_6180 (.Y(I6891),.A(g2962));
INVX1 NOT_6181 (.Y(g8292),.A(I13230));
INVX1 NOT_6182 (.Y(g2952),.A(g2455));
INVX1 NOT_6183 (.Y(I16956),.A(g11096));
INVX1 NOT_6184 (.Y(g3345),.A(I6531));
INVX1 NOT_6185 (.Y(I16376),.A(g10596));
INVX1 NOT_6186 (.Y(I13314),.A(g8260));
INVX1 NOT_6187 (.Y(g4284),.A(g3664));
INVX1 NOT_6188 (.Y(g7579),.A(I12053));
INVX1 NOT_6189 (.Y(g8526),.A(I13735));
INVX1 NOT_6190 (.Y(g10598),.A(I16273));
INVX1 NOT_6191 (.Y(g3763),.A(I6968));
INVX1 NOT_6192 (.Y(I10733),.A(g6099));
INVX1 NOT_6193 (.Y(g4545),.A(I7952));
INVX1 NOT_6194 (.Y(I11076),.A(g6649));
INVX1 NOT_6195 (.Y(I11085),.A(g6433));
INVX1 NOT_6196 (.Y(g3391),.A(g2896));
INVX1 NOT_6197 (.Y(g9733),.A(I14876));
INVX1 NOT_6198 (.Y(I15427),.A(g10088));
INVX1 NOT_6199 (.Y(I16095),.A(g10401));
INVX1 NOT_6200 (.Y(g4180),.A(I7357));
INVX1 NOT_6201 (.Y(g5490),.A(I8911));
INVX1 NOT_6202 (.Y(g9270),.A(I14485));
INVX1 NOT_6203 (.Y(g4380),.A(I7701));
INVX1 NOT_6204 (.Y(g11427),.A(I17334));
INVX1 NOT_6205 (.Y(g5166),.A(g4682));
INVX1 NOT_6206 (.Y(I11596),.A(g6831));
INVX1 NOT_6207 (.Y(g4591),.A(g3829));
INVX1 NOT_6208 (.Y(I15632),.A(g10184));
INVX1 NOT_6209 (.Y(g11366),.A(I17191));
INVX1 NOT_6210 (.Y(g3637),.A(I6818));
INVX1 NOT_6211 (.Y(I7216),.A(g2952));
INVX1 NOT_6212 (.Y(g7752),.A(I12421));
INVX1 NOT_6213 (.Y(g11632),.A(I17710));
INVX1 NOT_6214 (.Y(g8484),.A(g8336));
INVX1 NOT_6215 (.Y(I16181),.A(g10491));
INVX1 NOT_6216 (.Y(I10630),.A(g5889));
INVX1 NOT_6217 (.Y(g8439),.A(I13615));
INVX1 NOT_6218 (.Y(g2004),.A(I4820));
INVX1 NOT_6219 (.Y(I10693),.A(g6068));
INVX1 NOT_6220 (.Y(g6836),.A(I10888));
INVX1 NOT_6221 (.Y(I12372),.A(g7137));
INVX1 NOT_6222 (.Y(g7917),.A(g7497));
INVX1 NOT_6223 (.Y(g2986),.A(I6220));
INVX1 NOT_6224 (.Y(g3307),.A(I6480));
INVX1 NOT_6225 (.Y(g9473),.A(g9103));
INVX1 NOT_6226 (.Y(I7671),.A(g3351));
INVX1 NOT_6227 (.Y(g2647),.A(g1993));
INVX1 NOT_6228 (.Y(g10159),.A(I15473));
INVX1 NOT_6229 (.Y(g4420),.A(I7766));
INVX1 NOT_6230 (.Y(g10125),.A(I15377));
INVX1 NOT_6231 (.Y(g10532),.A(g10473));
INVX1 NOT_6232 (.Y(g10901),.A(g10802));
INVX1 NOT_6233 (.Y(I10009),.A(g5542));
INVX1 NOT_6234 (.Y(g5649),.A(I9108));
INVX1 NOT_6235 (.Y(g3359),.A(I6543));
INVX1 NOT_6236 (.Y(I15403),.A(g10069));
INVX1 NOT_6237 (.Y(g1965),.A(g119));
INVX1 NOT_6238 (.Y(g4507),.A(g3546));
INVX1 NOT_6239 (.Y(g5348),.A(I8815));
INVX1 NOT_6240 (.Y(g6967),.A(I11119));
INVX1 NOT_6241 (.Y(I5555),.A(g110));
INVX1 NOT_6242 (.Y(I11269),.A(g6545));
INVX1 NOT_6243 (.Y(g9980),.A(I15181));
INVX1 NOT_6244 (.Y(g2764),.A(I5850));
INVX1 NOT_6245 (.Y(I8462),.A(g4475));
INVX1 NOT_6246 (.Y(g11403),.A(I17252));
INVX1 NOT_6247 (.Y(g10158),.A(I15470));
INVX1 NOT_6248 (.Y(g11547),.A(g11519));
INVX1 NOT_6249 (.Y(g7042),.A(I11211));
INVX1 NOT_6250 (.Y(I11773),.A(g7257));
INVX1 NOT_6251 (.Y(g10783),.A(I16479));
INVX1 NOT_6252 (.Y(g4794),.A(I8164));
INVX1 NOT_6253 (.Y(I11942),.A(g6909));
INVX1 NOT_6254 (.Y(I13773),.A(g8384));
INVX1 NOT_6255 (.Y(I5792),.A(g2080));
INVX1 NOT_6256 (.Y(g7442),.A(g7237));
INVX1 NOT_6257 (.Y(g8702),.A(g8664));
INVX1 NOT_6258 (.Y(I13341),.A(g8210));
INVX1 NOT_6259 (.Y(I12790),.A(g7618));
INVX1 NOT_6260 (.Y(g7786),.A(I12523));
INVX1 NOT_6261 (.Y(g2503),.A(g1872));
INVX1 NOT_6262 (.Y(g3757),.A(I6952));
INVX1 NOT_6263 (.Y(I9352),.A(g4944));
INVX1 NOT_6264 (.Y(I17312),.A(g11392));
INVX1 NOT_6265 (.Y(g10353),.A(I15823));
INVX1 NOT_6266 (.Y(g3416),.A(g3144));
INVX1 NOT_6267 (.Y(g6993),.A(I11135));
INVX1 NOT_6268 (.Y(I11180),.A(g6506));
INVX1 NOT_6269 (.Y(I16190),.A(g10493));
INVX1 NOT_6270 (.Y(I14485),.A(g8883));
INVX1 NOT_6271 (.Y(g7364),.A(I11740));
INVX1 NOT_6272 (.Y(I6815),.A(g2755));
INVX1 NOT_6273 (.Y(I9717),.A(g5426));
INVX1 NOT_6274 (.Y(I15551),.A(g10080));
INVX1 NOT_6275 (.Y(I14555),.A(g9009));
INVX1 NOT_6276 (.Y(g3522),.A(g3164));
INVX1 NOT_6277 (.Y(g8952),.A(I14309));
INVX1 NOT_6278 (.Y(g11572),.A(g11561));
INVX1 NOT_6279 (.Y(I11734),.A(g7024));
INVX1 NOT_6280 (.Y(g8276),.A(I13200));
INVX1 NOT_6281 (.Y(g3811),.A(I7029));
INVX1 NOT_6282 (.Y(g2224),.A(g695));
INVX1 NOT_6283 (.Y(I6097),.A(g2391));
INVX1 NOT_6284 (.Y(g5063),.A(g4363));
INVX1 NOT_6285 (.Y(I10914),.A(g6728));
INVX1 NOT_6286 (.Y(g7454),.A(g7148));
INVX1 NOT_6287 (.Y(I6726),.A(g3306));
INVX1 NOT_6288 (.Y(I14570),.A(g9028));
INVX1 NOT_6289 (.Y(I9893),.A(g5557));
INVX1 NOT_6290 (.Y(I13335),.A(g8206));
INVX1 NOT_6291 (.Y(g7770),.A(I12475));
INVX1 NOT_6292 (.Y(I14914),.A(g9533));
INVX1 NOT_6293 (.Y(g4515),.A(I7916));
INVX1 NOT_6294 (.Y(g4204),.A(I7429));
INVX1 NOT_6295 (.Y(I15127),.A(g9919));
INVX1 NOT_6296 (.Y(I16546),.A(g10724));
INVX1 NOT_6297 (.Y(g8561),.A(I13776));
INVX1 NOT_6298 (.Y(g2320),.A(g18));
INVX1 NOT_6299 (.Y(I10907),.A(g6705));
INVX1 NOT_6300 (.Y(g7725),.A(I12360));
INVX1 NOT_6301 (.Y(I8842),.A(g4556));
INVX1 NOT_6302 (.Y(g7532),.A(I11932));
INVX1 NOT_6303 (.Y(I7308),.A(g3070));
INVX1 NOT_6304 (.Y(g3874),.A(g2920));
INVX1 NOT_6305 (.Y(I8192),.A(g3566));
INVX1 NOT_6306 (.Y(I12208),.A(g7124));
INVX1 NOT_6307 (.Y(I8298),.A(g4437));
INVX1 NOT_6308 (.Y(I8085),.A(g3664));
INVX1 NOT_6309 (.Y(I13965),.A(g8451));
INVX1 NOT_6310 (.Y(g8004),.A(I12838));
INVX1 NOT_6311 (.Y(g6921),.A(I11037));
INVX1 NOT_6312 (.Y(g8986),.A(I14379));
INVX1 NOT_6313 (.Y(I5494),.A(g1690));
INVX1 NOT_6314 (.Y(I13131),.A(g7979));
INVX1 NOT_6315 (.Y(I14239),.A(g8803));
INVX1 NOT_6316 (.Y(I15956),.A(g10402));
INVX1 NOT_6317 (.Y(g2617),.A(g1997));
INVX1 NOT_6318 (.Y(g2906),.A(I6071));
INVX1 NOT_6319 (.Y(I14567),.A(g9027));
INVX1 NOT_6320 (.Y(g2789),.A(g2276));
INVX1 NOT_6321 (.Y(g5619),.A(g4840));
INVX1 NOT_6322 (.Y(g5167),.A(g4682));
INVX1 NOT_6323 (.Y(I15980),.A(g10414));
AND2X1 AND2_0 (.Y(g11103),.A(g2250),.B(g10937));
AND2X1 AND2_1 (.Y(g9900),.A(g9845),.B(g8327));
AND2X1 AND2_2 (.Y(g11095),.A(g845),.B(g10950));
AND2X1 AND2_3 (.Y(g3880),.A(g3186),.B(g2023));
AND2X1 AND2_4 (.Y(g4973),.A(g1645),.B(g4467));
AND2X1 AND2_5 (.Y(g7389),.A(g7001),.B(g3880));
AND2X1 AND2_6 (.Y(g7888),.A(g7465),.B(g7025));
AND2X1 AND2_7 (.Y(g4969),.A(g1642),.B(g4463));
AND2X1 AND2_8 (.Y(g8224),.A(g1882),.B(g7887));
AND2X1 AND2_9 (.Y(g2892),.A(g1980),.B(g1976));
AND2X1 AND2_10 (.Y(g5686),.A(g158),.B(g5361));
AND2X1 AND2_11 (.Y(g10308),.A(g10217),.B(g9085));
AND2X1 AND2_12 (.Y(g4123),.A(g2695),.B(g3037));
AND2X1 AND2_13 (.Y(g8120),.A(g1909),.B(g7944));
AND2X1 AND2_14 (.Y(g6788),.A(g287),.B(g5876));
AND2X1 AND2_15 (.Y(g5598),.A(g778),.B(g4824));
AND2X1 AND2_16 (.Y(g9694),.A(g278),.B(g9432));
AND2X1 AND2_17 (.Y(g10495),.A(g10431),.B(g3971));
AND2X1 AND2_18 (.Y(g2945),.A(g2411),.B(g1684));
AND2X1 AND2_19 (.Y(g11190),.A(g5623),.B(g11065));
AND2X1 AND2_20 (.Y(g8789),.A(g8639),.B(g8719));
AND2X1 AND2_21 (.Y(g9852),.A(g9728),.B(g9563));
AND2X1 AND2_22 (.Y(g5625),.A(g1053),.B(g4399));
AND2X1 AND2_23 (.Y(g4875),.A(g995),.B(g3914));
AND2X1 AND2_24 (.Y(g9701),.A(g1574),.B(g9474));
AND2X1 AND2_25 (.Y(g7138),.A(g6055),.B(g6707));
AND2X1 AND2_26 (.Y(g10752),.A(g10692),.B(g3586));
AND2X1 AND2_27 (.Y(g11211),.A(g11058),.B(g5534));
AND2X1 AND2_28 (.Y(g11024),.A(g435),.B(g10974));
AND2X1 AND2_29 (.Y(g8547),.A(g8307),.B(g7693));
AND2X1 AND2_30 (.Y(g10669),.A(g10577),.B(g9429));
AND2X1 AND2_31 (.Y(g7707),.A(g691),.B(g7206));
AND2X1 AND2_32 (.Y(g4884),.A(g3813),.B(g2971));
AND2X1 AND2_33 (.Y(g4839),.A(g225),.B(g3946));
AND2X1 AND2_34 (.Y(g9870),.A(g1561),.B(g9816));
AND2X1 AND2_35 (.Y(g6640),.A(g5281),.B(g5801));
AND2X1 AND2_36 (.Y(g9650),.A(g2797),.B(g9240));
AND2X1 AND2_37 (.Y(g5687),.A(g139),.B(g5361));
AND2X1 AND2_38 (.Y(g7957),.A(g2885),.B(g7527));
AND2X1 AND2_39 (.Y(g3512),.A(g2050),.B(g2971));
AND2X1 AND2_40 (.Y(g8244),.A(g7847),.B(g4336));
AND2X1 AND2_41 (.Y(g7449),.A(g6868),.B(g4355));
AND2X1 AND2_42 (.Y(g4235),.A(g1011),.B(g3914));
AND2X1 AND2_43 (.Y(g4343),.A(g345),.B(g3586));
AND2X1 AND2_44 (.Y(g11296),.A(g5482),.B(g11241));
AND2X1 AND2_45 (.Y(g9594),.A(g1),.B(g9292));
AND2X1 AND2_46 (.Y(g6829),.A(g213),.B(g6596));
AND2X1 AND2_47 (.Y(g4334),.A(g1160),.B(g3703));
AND2X1 AND2_48 (.Y(g9943),.A(g9923),.B(g9367));
AND2X1 AND2_49 (.Y(g5525),.A(g1721),.B(g4292));
AND2X1 AND2_50 (.Y(g4548),.A(g440),.B(g3990));
AND2X1 AND_tmp1 (.Y(ttmp1),.A(g6764),.B(g8858));
AND2X1 AND_tmp2 (.Y(g8876),.A(g8105),.B(ttmp1));
AND2X1 AND2_51 (.Y(g6733),.A(g5678),.B(g4324));
AND2X1 AND2_52 (.Y(g4804),.A(g476),.B(g3458));
AND2X1 AND2_53 (.Y(g10705),.A(g10564),.B(g4840));
AND2X1 AND2_54 (.Y(g9934),.A(g9913),.B(g9624));
AND2X1 AND2_55 (.Y(g6225),.A(g566),.B(g5082));
AND2X1 AND2_56 (.Y(g6324),.A(g1240),.B(g5949));
AND2X1 AND2_57 (.Y(g10686),.A(g10612),.B(g3863));
AND2X1 AND2_58 (.Y(g6540),.A(g1223),.B(g6072));
AND2X1 AND2_59 (.Y(g8663),.A(g8538),.B(g4013));
AND2X1 AND2_60 (.Y(g11581),.A(g1308),.B(g11539));
AND2X1 AND2_61 (.Y(g6206),.A(g560),.B(g5068));
AND2X1 AND2_62 (.Y(g4518),.A(g452),.B(g3975));
AND2X1 AND2_63 (.Y(g3989),.A(g248),.B(g3164));
AND2X1 AND2_64 (.Y(g7730),.A(g7260),.B(g2347));
AND2X1 AND2_65 (.Y(g5174),.A(g1235),.B(g4681));
AND2X1 AND2_66 (.Y(g7504),.A(g7148),.B(g2847));
AND2X1 AND2_67 (.Y(g7185),.A(g1887),.B(g6724));
AND2X1 AND2_68 (.Y(g2563),.A(I5689),.B(I5690));
AND2X1 AND2_69 (.Y(g7881),.A(g7612),.B(g3810));
AND2X1 AND2_70 (.Y(g11070),.A(g2008),.B(g10913));
AND2X1 AND2_71 (.Y(g9859),.A(g9736),.B(g9573));
AND2X1 AND_tmp3 (.Y(ttmp3),.A(g6764),.B(g8858));
AND2X1 AND_tmp4 (.Y(g8877),.A(g8103),.B(ttmp3));
AND2X1 AND2_72 (.Y(g11590),.A(g2274),.B(g11561));
AND2X1 AND2_73 (.Y(g6199),.A(g557),.B(g5062));
AND2X1 AND2_74 (.Y(g9266),.A(g8932),.B(g3398));
AND2X1 AND2_75 (.Y(g5545),.A(g1730),.B(g4321));
AND2X1 AND2_76 (.Y(g5180),.A(g4541),.B(g4533));
AND2X1 AND2_77 (.Y(g5591),.A(g1615),.B(g4514));
AND2X1 AND2_78 (.Y(g8556),.A(g8412),.B(g8029));
AND2X1 AND2_79 (.Y(g11094),.A(g374),.B(g10883));
AND2X1 AND2_80 (.Y(g5853),.A(g5044),.B(g1927));
AND2X1 AND2_81 (.Y(g6245),.A(g575),.B(g5098));
AND2X1 AND2_82 (.Y(g4360),.A(g1861),.B(g3748));
AND2X1 AND_tmp5 (.Y(ttmp5),.A(g6368),.B(g8828));
AND2X1 AND_tmp6 (.Y(g8930),.A(g8100),.B(ttmp5));
AND2X1 AND2_83 (.Y(g5507),.A(g4310),.B(g3528));
AND2X1 AND2_84 (.Y(g11150),.A(g3087),.B(g10913));
AND2X1 AND2_85 (.Y(g8464),.A(g8302),.B(g7416));
AND2X1 AND2_86 (.Y(g9692),.A(g272),.B(g9432));
AND2X1 AND2_87 (.Y(g4996),.A(g1428),.B(g4682));
AND2X1 AND2_88 (.Y(g7131),.A(g6044),.B(g6700));
AND2X1 AND2_89 (.Y(g11019),.A(g421),.B(g10974));
AND2X1 AND2_90 (.Y(g9960),.A(g9951),.B(g9536));
AND2X1 AND2_91 (.Y(g11196),.A(g4912),.B(g11068));
AND2X1 AND2_92 (.Y(g11018),.A(g7286),.B(g10974));
AND2X1 AND2_93 (.Y(g6819),.A(g243),.B(g6596));
AND2X1 AND2_94 (.Y(g10595),.A(g10550),.B(g4347));
AND2X1 AND2_95 (.Y(g10494),.A(g10433),.B(g3945));
AND2X1 AND2_96 (.Y(g10623),.A(g10544),.B(g4536));
AND2X1 AND2_97 (.Y(g4878),.A(g1868),.B(g3531));
AND2X1 AND2_98 (.Y(g5204),.A(g4838),.B(g2126));
AND2X1 AND2_99 (.Y(g8844),.A(g8609),.B(g8709));
AND2X1 AND2_100 (.Y(g6701),.A(g6185),.B(g4228));
AND2X1 AND2_101 (.Y(g10782),.A(g10725),.B(g5146));
AND2X1 AND2_102 (.Y(g5100),.A(g1791),.B(g4606));
AND2X1 AND2_103 (.Y(g4882),.A(g1089),.B(g3638));
AND2X1 AND2_104 (.Y(g8731),.A(g8622),.B(g7918));
AND2X1 AND2_105 (.Y(g6215),.A(g1504),.B(g5128));
AND2X1 AND2_106 (.Y(g6886),.A(g1932),.B(g6420));
AND2X1 AND2_107 (.Y(g3586),.A(g3323),.B(g2191));
AND2X1 AND2_108 (.Y(g8557),.A(g8415),.B(g8033));
AND2X1 AND_tmp7 (.Y(ttmp7),.A(g6778),.B(g8849));
AND2X1 AND_tmp8 (.Y(g8966),.A(g8081),.B(ttmp7));
AND2X1 AND2_109 (.Y(g8071),.A(g691),.B(g7826));
AND2X1 AND2_110 (.Y(g11597),.A(g11576),.B(g5446));
AND2X1 AND2_111 (.Y(g9828),.A(g9722),.B(g9785));
AND2X1 AND2_112 (.Y(g2918),.A(g2411),.B(g1672));
AND2X1 AND2_113 (.Y(g9830),.A(g9725),.B(g9785));
AND2X1 AND_tmp9 (.Y(ttmp9),.A(g6368),.B(g8828));
AND2X1 AND_tmp10 (.Y(g8955),.A(g8110),.B(ttmp9));
AND2X1 AND2_114 (.Y(g9592),.A(g4),.B(g9292));
AND2X1 AND2_115 (.Y(g5123),.A(g1618),.B(g4669));
AND2X1 AND2_116 (.Y(g7059),.A(g6078),.B(g6714));
AND2X1 AND2_117 (.Y(g8254),.A(g2773),.B(g7909));
AND2X1 AND2_118 (.Y(g7459),.A(g7148),.B(g2814));
AND2X1 AND2_119 (.Y(g11102),.A(g861),.B(g10950));
AND2X1 AND2_120 (.Y(g7718),.A(g709),.B(g7221));
AND2X1 AND2_121 (.Y(g7535),.A(g7148),.B(g2874));
AND2X1 AND2_122 (.Y(g9703),.A(g1577),.B(g9474));
AND2X1 AND2_123 (.Y(g5528),.A(g4322),.B(g3537));
AND2X1 AND2_124 (.Y(g5151),.A(g4478),.B(g2733));
AND2X1 AND2_125 (.Y(g9932),.A(g9911),.B(g9624));
AND2X1 AND2_126 (.Y(g5530),.A(g1636),.B(g4305));
AND2X1 AND2_127 (.Y(g3506),.A(g986),.B(g2760));
AND2X1 AND2_128 (.Y(g8769),.A(g8629),.B(g5151));
AND2X1 AND2_129 (.Y(g6887),.A(g6187),.B(g6566));
AND2X1 AND2_130 (.Y(g6228),.A(g5605),.B(g713));
AND2X1 AND2_131 (.Y(g6322),.A(g1275),.B(g5949));
AND2X1 AND2_132 (.Y(g3111),.A(I6337),.B(I6338));
AND2X1 AND_tmp11 (.Y(ttmp11),.A(g6778),.B(g8849));
AND2X1 AND_tmp12 (.Y(g8967),.A(g8085),.B(ttmp11));
AND2X1 AND2_133 (.Y(g5010),.A(g1458),.B(g4640));
AND2X1 AND2_134 (.Y(g3275),.A(g115),.B(g2356));
AND2X1 AND2_135 (.Y(g10809),.A(g4811),.B(g10754));
AND2X1 AND2_136 (.Y(g2895),.A(g2411),.B(g1678));
AND2X1 AND2_137 (.Y(g7721),.A(g736),.B(g7237));
AND2X1 AND2_138 (.Y(g9866),.A(g1549),.B(g9802));
AND2X1 AND2_139 (.Y(g9716),.A(g1534),.B(g9490));
AND2X1 AND2_140 (.Y(g10808),.A(g10744),.B(g3829));
AND2X1 AND2_141 (.Y(g3374),.A(g1231),.B(g3047));
AND2X1 AND2_142 (.Y(g4492),.A(g1786),.B(g3685));
AND2X1 AND2_143 (.Y(g8822),.A(g8614),.B(g8752));
AND2X1 AND2_144 (.Y(g10560),.A(g10487),.B(g4575));
AND2X1 AND_tmp13 (.Y(ttmp13),.A(g3517),.B(g11422));
AND2X1 AND_tmp14 (.Y(g11456),.A(g3765),.B(ttmp13));
AND2X1 AND2_145 (.Y(g9848),.A(g9724),.B(g9557));
AND2X1 AND2_146 (.Y(g4714),.A(g646),.B(g3333));
AND2X1 AND2_147 (.Y(g6550),.A(g1231),.B(g6089));
AND2X1 AND2_148 (.Y(g5172),.A(g4555),.B(g4549));
AND2X1 AND2_149 (.Y(g10642),.A(g10612),.B(g3829));
AND2X1 AND2_150 (.Y(g3284),.A(g2531),.B(g677));
AND2X1 AND2_151 (.Y(g9699),.A(g284),.B(g9432));
AND2X1 AND2_152 (.Y(g9855),.A(g302),.B(g9772));
AND2X1 AND2_153 (.Y(g5618),.A(g1630),.B(g4551));
AND2X1 AND2_154 (.Y(g6891),.A(g1950),.B(g6435));
AND2X1 AND2_155 (.Y(g7940),.A(g7620),.B(g4013));
AND2X1 AND2_156 (.Y(g11085),.A(g312),.B(g10897));
AND2X1 AND2_157 (.Y(g4736),.A(g396),.B(g3379));
AND2X1 AND2_158 (.Y(g4968),.A(g1432),.B(g4682));
AND2X1 AND2_159 (.Y(g8837),.A(g8646),.B(g8697));
AND2X1 AND2_160 (.Y(g9644),.A(g1182),.B(g9125));
AND2X1 AND2_161 (.Y(g5804),.A(g1546),.B(g5261));
AND2X1 AND2_162 (.Y(g8462),.A(g8300),.B(g7406));
AND2X1 AND_tmp15 (.Y(ttmp15),.A(g2562),.B(g2570));
AND2X1 AND_tmp16 (.Y(ttmp16),.A(g2549),.B(ttmp15));
AND2X1 AND_tmp17 (.Y(I6330),.A(g2556),.B(ttmp16));
AND2X1 AND2_163 (.Y(g11156),.A(g333),.B(g10934));
AND2X1 AND2_164 (.Y(g6342),.A(g293),.B(g5886));
AND2X1 AND2_165 (.Y(g9867),.A(g1552),.B(g9807));
AND2X1 AND2_166 (.Y(g9717),.A(g1537),.B(g9490));
AND2X1 AND2_167 (.Y(g4871),.A(g1864),.B(g3523));
AND2X1 AND2_168 (.Y(g10454),.A(g10435),.B(g3411));
AND2X1 AND2_169 (.Y(g4722),.A(g426),.B(g3353));
AND2X1 AND2_170 (.Y(g7741),.A(g6961),.B(g3880));
AND2X1 AND2_171 (.Y(g4500),.A(g1357),.B(g3941));
AND2X1 AND2_172 (.Y(g9386),.A(g1327),.B(g9151));
AND2X1 AND2_173 (.Y(g8842),.A(g8607),.B(g8707));
AND2X1 AND2_174 (.Y(g9599),.A(g8),.B(g9292));
AND2X1 AND2_175 (.Y(g9274),.A(g8974),.B(g5708));
AND2X1 AND2_176 (.Y(g5518),.A(g4317),.B(g3532));
AND2X1 AND2_177 (.Y(g9614),.A(g1197),.B(g9111));
AND2X1 AND2_178 (.Y(g4838),.A(g3275),.B(g4122));
AND2X1 AND2_179 (.Y(g9125),.A(g8966),.B(g6674));
AND2X1 AND2_180 (.Y(g7217),.A(g4610),.B(g6432));
AND2X1 AND2_181 (.Y(g11557),.A(g2707),.B(g11519));
AND2X1 AND2_182 (.Y(g2911),.A(g2411),.B(g1675));
AND2X1 AND2_183 (.Y(g11210),.A(g11078),.B(g4515));
AND2X1 AND2_184 (.Y(g7466),.A(g7148),.B(g2821));
AND2X1 AND2_185 (.Y(g9939),.A(g9918),.B(g9367));
AND2X1 AND2_186 (.Y(g11279),.A(g4939),.B(g11200));
AND2X1 AND_tmp18 (.Y(ttmp18),.A(g10440),.B(I16145));
AND2X1 AND_tmp19 (.Y(g10518),.A(g10513),.B(ttmp18));
AND2X1 AND2_187 (.Y(g4477),.A(g1129),.B(g3878));
AND2X1 AND2_188 (.Y(g8708),.A(g7605),.B(g8592));
AND2X1 AND2_189 (.Y(g7055),.A(g5900),.B(g6579));
AND2X1 AND2_190 (.Y(g5264),.A(g1095),.B(g4763));
AND2X1 AND2_191 (.Y(g6329),.A(g1265),.B(g5949));
AND2X1 AND2_192 (.Y(g6828),.A(g1377),.B(g6596));
AND2X1 AND2_193 (.Y(g8176),.A(g5299),.B(g7853));
AND2X1 AND2_194 (.Y(g6830),.A(g1380),.B(g6596));
AND2X1 AND2_195 (.Y(g8005),.A(g7510),.B(g6871));
AND2X1 AND2_196 (.Y(g4099),.A(g770),.B(g3281));
AND2X1 AND2_197 (.Y(g11601),.A(g1351),.B(g11574));
AND2X1 AND2_198 (.Y(g11187),.A(g5597),.B(g11061));
AND2X1 AND2_199 (.Y(g6746),.A(g6228),.B(g6166));
AND2X1 AND2_200 (.Y(g6221),.A(g782),.B(g5598));
AND2X1 AND2_201 (.Y(g8765),.A(g8630),.B(g5151));
AND2X1 AND2_202 (.Y(g9622),.A(g1200),.B(g9111));
AND2X1 AND2_203 (.Y(g11143),.A(g10923),.B(g4567));
AND2X1 AND2_204 (.Y(g9904),.A(g9886),.B(g9676));
AND2X1 AND2_205 (.Y(g8733),.A(g8625),.B(g7920));
AND2X1 AND_tmp20 (.Y(ttmp20),.A(g6368),.B(g8858));
AND2X1 AND_tmp21 (.Y(g8974),.A(g8094),.B(ttmp20));
AND2X1 AND2_206 (.Y(g6624),.A(g348),.B(g6171));
AND2X1 AND2_207 (.Y(g11169),.A(g530),.B(g11112));
AND2X1 AND2_208 (.Y(g8073),.A(g709),.B(g7826));
AND2X1 AND2_209 (.Y(g9841),.A(g9706),.B(g9512));
AND2X1 AND2_210 (.Y(g5882),.A(g5592),.B(g3829));
AND2X1 AND2_211 (.Y(g8796),.A(g8645),.B(g8725));
AND2X1 AND2_212 (.Y(g11168),.A(g534),.B(g11112));
AND2X1 AND2_213 (.Y(g4269),.A(g1015),.B(g3914));
AND2X1 AND2_214 (.Y(g5271),.A(g727),.B(g4772));
AND2X1 AND2_215 (.Y(g10348),.A(g10272),.B(g3705));
AND2X1 AND2_216 (.Y(g5611),.A(g1047),.B(g4382));
AND2X1 AND2_217 (.Y(g8069),.A(g673),.B(g7826));
AND2X1 AND2_218 (.Y(g9695),.A(g1567),.B(g9474));
AND2X1 AND2_219 (.Y(g10304),.A(g10211),.B(g9079));
AND2X1 AND2_220 (.Y(g8469),.A(g8305),.B(g7422));
AND2X1 AND2_221 (.Y(g4712),.A(g1071),.B(g3638));
AND2X1 AND2_222 (.Y(g6576),.A(g5762),.B(g5503));
AND2X1 AND2_223 (.Y(g10622),.A(g10543),.B(g4525));
AND2X1 AND2_224 (.Y(g11015),.A(g5217),.B(g10827));
AND2X1 AND2_225 (.Y(g5674),.A(g148),.B(g5361));
AND2X1 AND2_226 (.Y(g9359),.A(g1308),.B(g9173));
AND2X1 AND2_227 (.Y(g9223),.A(g6454),.B(g8960));
AND2X1 AND2_228 (.Y(g11556),.A(g2701),.B(g11519));
AND2X1 AND2_229 (.Y(g9858),.A(g1595),.B(g9774));
AND2X1 AND2_230 (.Y(g5541),.A(g4331),.B(g3582));
AND2X1 AND2_231 (.Y(g4534),.A(g363),.B(g3586));
AND2X1 AND2_232 (.Y(g6198),.A(g1499),.B(g5128));
AND2X1 AND2_233 (.Y(g6747),.A(g2214),.B(g5897));
AND2X1 AND2_234 (.Y(g6699),.A(g6177),.B(g4221));
AND2X1 AND2_235 (.Y(g6855),.A(g1964),.B(g6392));
AND2X1 AND2_236 (.Y(g3804),.A(g3098),.B(g2203));
AND2X1 AND2_237 (.Y(g5680),.A(g153),.B(g5361));
AND2X1 AND2_238 (.Y(g9642),.A(g2654),.B(g9240));
AND2X1 AND2_239 (.Y(g5744),.A(g1528),.B(g5191));
AND2X1 AND2_240 (.Y(g10333),.A(g10262),.B(g3307));
AND2X1 AND2_241 (.Y(g8399),.A(g6094),.B(g8229));
AND2X1 AND2_242 (.Y(g9447),.A(g1762),.B(g9030));
AND2X1 AND2_243 (.Y(g4903),.A(g1849),.B(g4243));
AND2X1 AND2_244 (.Y(g11178),.A(g516),.B(g11112));
AND2X1 AND2_245 (.Y(g8510),.A(g8414),.B(g7972));
AND2X1 AND2_246 (.Y(g8245),.A(g7850),.B(g4339));
AND2X1 AND2_247 (.Y(g6319),.A(g1296),.B(g5949));
AND2X1 AND2_248 (.Y(g11186),.A(g5594),.B(g11059));
AND2X1 AND2_249 (.Y(g3908),.A(g186),.B(g3164));
AND2X1 AND2_250 (.Y(g2951),.A(g2411),.B(g1681));
AND2X1 AND2_251 (.Y(g6352),.A(g278),.B(g5894));
AND2X1 AND2_252 (.Y(g9595),.A(g901),.B(g9205));
AND2X1 AND2_253 (.Y(g4831),.A(g810),.B(g4109));
AND2X1 AND2_254 (.Y(g5492),.A(g1654),.B(g4263));
AND2X1 AND2_255 (.Y(g9272),.A(g8934),.B(g3424));
AND2X1 AND2_256 (.Y(g10312),.A(g10220),.B(g9094));
AND2X1 AND2_257 (.Y(g6186),.A(g546),.B(g5042));
AND2X1 AND2_258 (.Y(g9612),.A(g2652),.B(g9240));
AND2X1 AND2_259 (.Y(g9417),.A(g1738),.B(g9052));
AND2X1 AND2_260 (.Y(g9935),.A(g9914),.B(g9624));
AND2X1 AND2_261 (.Y(g8701),.A(g7597),.B(g8582));
AND2X1 AND2_262 (.Y(g10745),.A(g10658),.B(g3586));
AND2X1 AND2_263 (.Y(g11216),.A(g956),.B(g11162));
AND2X1 AND2_264 (.Y(g9328),.A(g8971),.B(g5708));
AND2X1 AND2_265 (.Y(g11587),.A(g1327),.B(g11546));
AND2X1 AND2_266 (.Y(g6821),.A(g237),.B(g6596));
AND2X1 AND2_267 (.Y(g6325),.A(g1245),.B(g5949));
AND2X1 AND2_268 (.Y(g4560),.A(g431),.B(g4002));
AND2X1 AND2_269 (.Y(g7368),.A(g6980),.B(g3880));
AND2X1 AND2_270 (.Y(g6083),.A(g552),.B(g5619));
AND2X1 AND2_271 (.Y(g6544),.A(g1227),.B(g6081));
AND2X1 AND2_272 (.Y(g5476),.A(g1615),.B(g4237));
AND2X1 AND2_273 (.Y(g7743),.A(g6967),.B(g3880));
AND2X1 AND2_274 (.Y(g4869),.A(g1083),.B(g3638));
AND2X1 AND2_275 (.Y(g5722),.A(g1598),.B(g5144));
AND2X1 AND2_276 (.Y(g6790),.A(g5813),.B(g4398));
AND2X1 AND2_277 (.Y(g8408),.A(g704),.B(g8139));
AND2X1 AND2_278 (.Y(g10761),.A(g10700),.B(g10699));
AND2X1 AND2_279 (.Y(g7734),.A(g6944),.B(g3880));
AND2X1 AND2_280 (.Y(g8136),.A(g7926),.B(g7045));
AND2X1 AND2_281 (.Y(g6187),.A(g5569),.B(g2340));
AND2X1 AND2_282 (.Y(g4752),.A(g401),.B(g3385));
AND2X1 AND2_283 (.Y(g9902),.A(g9894),.B(g9392));
AND2X1 AND2_284 (.Y(g8768),.A(g8623),.B(g5151));
AND2X1 AND2_285 (.Y(g5500),.A(g1657),.B(g4272));
AND2X1 AND2_286 (.Y(g2496),.A(g374),.B(g369));
AND2X1 AND2_287 (.Y(g6756),.A(g3010),.B(g5877));
AND2X1 AND_tmp22 (.Y(ttmp22),.A(g6764),.B(g8858));
AND2X1 AND_tmp23 (.Y(g8972),.A(g8085),.B(ttmp22));
AND2X1 AND2_288 (.Y(g6622),.A(g336),.B(g6165));
AND2X1 AND2_289 (.Y(g11639),.A(g11612),.B(g7897));
AND2X1 AND2_290 (.Y(g9366),.A(g1311),.B(g9173));
AND2X1 AND2_291 (.Y(g11230),.A(g471),.B(g11062));
AND2X1 AND2_292 (.Y(g10328),.A(g10252),.B(g3307));
AND2X1 AND2_293 (.Y(g5024),.A(g1284),.B(g4513));
AND2X1 AND2_294 (.Y(g4364),.A(g1215),.B(g3756));
AND2X1 AND2_295 (.Y(g9649),.A(g916),.B(g9205));
AND2X1 AND2_296 (.Y(g5795),.A(g1543),.B(g5251));
AND2X1 AND2_297 (.Y(g5737),.A(g1524),.B(g5183));
AND2X1 AND2_298 (.Y(g6841),.A(g1400),.B(g6596));
AND2X1 AND2_299 (.Y(g4054),.A(g1753),.B(g2793));
AND2X1 AND2_300 (.Y(g6345),.A(g5823),.B(g4426));
AND2X1 AND2_301 (.Y(g11391),.A(g11275),.B(g7912));
AND2X1 AND2_302 (.Y(g9851),.A(g296),.B(g9770));
AND2X1 AND2_303 (.Y(g6763),.A(g5802),.B(g4381));
AND2X1 AND2_304 (.Y(g4770),.A(g416),.B(g3415));
AND2X1 AND_tmp24 (.Y(ttmp24),.A(g10509),.B(g10507));
AND2X1 AND_tmp25 (.Y(I16142),.A(g10511),.B(ttmp24));
AND2X1 AND2_305 (.Y(g9698),.A(g1571),.B(g9474));
AND2X1 AND2_306 (.Y(g4725),.A(g1032),.B(g3914));
AND2X1 AND2_307 (.Y(g5477),.A(g1887),.B(g4241));
AND2X1 AND2_308 (.Y(g9964),.A(g9954),.B(g9536));
AND2X1 AND2_309 (.Y(g5523),.A(g1663),.B(g4290));
AND2X1 AND2_310 (.Y(g4553),.A(g435),.B(g3995));
AND2X1 AND2_311 (.Y(g8550),.A(g8402),.B(g8011));
AND2X1 AND2_312 (.Y(g8845),.A(g8611),.B(g8711));
AND2X1 AND2_313 (.Y(g2081),.A(g932),.B(g928));
AND2X1 AND2_314 (.Y(g6359),.A(g281),.B(g5898));
AND2X1 AND2_315 (.Y(g11586),.A(g1324),.B(g11545));
AND2X1 AND2_316 (.Y(g11007),.A(g5147),.B(g10827));
AND2X1 AND2_317 (.Y(g5104),.A(g1796),.B(g4608));
AND2X1 AND2_318 (.Y(g5099),.A(g4821),.B(g3829));
AND2X1 AND2_319 (.Y(g6757),.A(g2221),.B(g5919));
AND2X1 AND2_320 (.Y(g5499),.A(g1627),.B(g4270));
AND2X1 AND2_321 (.Y(g4389),.A(g3529),.B(g3092));
AND2X1 AND2_322 (.Y(g6416),.A(g3497),.B(g5774));
AND2X1 AND2_323 (.Y(g9720),.A(g1546),.B(g9490));
AND2X1 AND2_324 (.Y(g4990),.A(g1444),.B(g4682));
AND2X1 AND2_325 (.Y(g9619),.A(g2772),.B(g9010));
AND2X1 AND_tmp26 (.Y(ttmp26),.A(g2689),.B(g2701));
AND2X1 AND_tmp27 (.Y(ttmp27),.A(g2677),.B(ttmp26));
AND2X1 AND_tmp28 (.Y(I6630),.A(g2683),.B(ttmp27));
AND2X1 AND2_326 (.Y(g6047),.A(g2017),.B(g4977));
AND2X1 AND2_327 (.Y(g9652),.A(g953),.B(g9223));
AND2X1 AND_tmp29 (.Y(ttmp29),.A(g10469),.B(I16142));
AND2X1 AND_tmp30 (.Y(g10515),.A(g10505),.B(ttmp29));
AND2X1 AND2_328 (.Y(g9843),.A(g9711),.B(g9519));
AND2X1 AND2_329 (.Y(g5273),.A(g1074),.B(g4776));
AND2X1 AND2_330 (.Y(g11465),.A(g11434),.B(g5446));
AND2X1 AND2_331 (.Y(g5044),.A(g4348),.B(g1918));
AND2X1 AND2_332 (.Y(g11237),.A(g5472),.B(g11109));
AND2X1 AND2_333 (.Y(g9834),.A(g9731),.B(g9785));
AND2X1 AND2_334 (.Y(g6654),.A(g363),.B(g6214));
AND2X1 AND2_335 (.Y(g5444),.A(g1041),.B(g4880));
AND2X1 AND2_336 (.Y(g3714),.A(g1690),.B(g2991));
AND2X1 AND2_337 (.Y(g11340),.A(g11285),.B(g4424));
AND2X1 AND2_338 (.Y(g9598),.A(g2086),.B(g9274));
AND2X1 AND2_339 (.Y(g8097),.A(g6200),.B(g7851));
AND2X1 AND2_340 (.Y(g8726),.A(g8608),.B(g7913));
AND2X1 AND2_341 (.Y(g6880),.A(g4816),.B(g6562));
AND2X1 AND2_342 (.Y(g4338),.A(g1157),.B(g3707));
AND2X1 AND2_343 (.Y(g5543),.A(g4874),.B(g4312));
AND2X1 AND_tmp31 (.Y(ttmp31),.A(g6368),.B(g8828));
AND2X1 AND_tmp32 (.Y(g8960),.A(g8085),.B(ttmp31));
AND2X1 AND2_344 (.Y(g4109),.A(g806),.B(g3287));
AND2X1 AND2_345 (.Y(g10759),.A(g10698),.B(g10697));
AND2X1 AND2_346 (.Y(g9938),.A(g9917),.B(g9367));
AND2X1 AND2_347 (.Y(g10758),.A(g10652),.B(g4013));
AND2X1 AND2_348 (.Y(g4759),.A(g406),.B(g3392));
AND2X1 AND2_349 (.Y(g9909),.A(g9891),.B(g9804));
AND2X1 AND2_350 (.Y(g7127),.A(g6663),.B(g2241));
AND2X1 AND2_351 (.Y(g11165),.A(g476),.B(g11112));
AND2X1 AND2_352 (.Y(g6234),.A(g2244),.B(g5151));
AND2X1 AND2_353 (.Y(g6328),.A(g1260),.B(g5949));
AND2X1 AND2_354 (.Y(g8401),.A(g677),.B(g8124));
AND2X1 AND2_355 (.Y(g11006),.A(g5125),.B(g10827));
AND2X1 AND2_356 (.Y(g4865),.A(g1080),.B(g3638));
AND2X1 AND2_357 (.Y(g4715),.A(g1077),.B(g3638));
AND2X1 AND_tmp33 (.Y(ttmp33),.A(g3753),.B(g2325));
AND2X1 AND_tmp34 (.Y(g4604),.A(g3056),.B(ttmp33));
AND2X1 AND2_358 (.Y(g5513),.A(g1675),.B(g4282));
AND2X1 AND2_359 (.Y(g11222),.A(g965),.B(g11055));
AND2X1 AND2_360 (.Y(g4498),.A(g1145),.B(g3940));
AND2X1 AND2_361 (.Y(g6554),.A(g5075),.B(g6183));
AND2X1 AND2_362 (.Y(g7732),.A(g6935),.B(g3880));
AND2X1 AND2_363 (.Y(g9586),.A(g2727),.B(g9173));
AND2X1 AND_tmp35 (.Y(ttmp35),.A(g4401),.B(g4104));
AND2X1 AND_tmp36 (.Y(g5178),.A(g2047),.B(ttmp35));
AND2X1 AND2_364 (.Y(g4584),.A(g3710),.B(g2322));
AND2X1 AND2_365 (.Y(g7472),.A(g7148),.B(g2829));
AND2X1 AND2_366 (.Y(g11253),.A(g981),.B(g11072));
AND2X1 AND2_367 (.Y(g5182),.A(g1240),.B(g4713));
AND2X1 AND2_368 (.Y(g9860),.A(g1598),.B(g9775));
AND2X1 AND2_369 (.Y(g8703),.A(g7601),.B(g8585));
AND2X1 AND2_370 (.Y(g11600),.A(g1346),.B(g11573));
AND2X1 AND2_371 (.Y(g9710),.A(g1586),.B(g9474));
AND2X1 AND2_372 (.Y(g9645),.A(g1203),.B(g9111));
AND2X1 AND2_373 (.Y(g11236),.A(g5469),.B(g11108));
AND2X1 AND2_374 (.Y(g4162),.A(g3106),.B(g2971));
AND2X1 AND2_375 (.Y(g6090),.A(g553),.B(g5627));
AND2X1 AND2_376 (.Y(g9691),.A(g269),.B(g9432));
AND2X1 AND2_377 (.Y(g11372),.A(g11316),.B(g4266));
AND2X1 AND2_378 (.Y(g6823),.A(g1368),.B(g6596));
AND2X1 AND2_379 (.Y(g11175),.A(g501),.B(g11112));
AND2X1 AND2_380 (.Y(g8068),.A(g664),.B(g7826));
AND2X1 AND2_381 (.Y(g9607),.A(g12),.B(g9274));
AND2X1 AND2_382 (.Y(g9962),.A(g9952),.B(g9536));
AND2X1 AND2_383 (.Y(g6348),.A(g296),.B(g5891));
AND2X1 AND2_384 (.Y(g9659),.A(g956),.B(g9223));
AND2X1 AND2_385 (.Y(g9358),.A(g1318),.B(g9151));
AND2X1 AND2_386 (.Y(g3104),.A(I6316),.B(I6317));
AND2X1 AND2_387 (.Y(g4486),.A(g1711),.B(g3910));
AND2X1 AND2_388 (.Y(g9587),.A(g892),.B(g8995));
AND2X1 AND2_389 (.Y(g5632),.A(g1636),.B(g4563));
AND2X1 AND2_390 (.Y(g9111),.A(g8965),.B(g6674));
AND2X1 AND2_391 (.Y(g4881),.A(g991),.B(g3914));
AND2X1 AND2_392 (.Y(g11209),.A(g11074),.B(g9448));
AND2X1 AND2_393 (.Y(g8848),.A(g8715),.B(g8713));
AND2X1 AND2_394 (.Y(g4070),.A(g3263),.B(g2330));
AND2X1 AND2_395 (.Y(g6463),.A(g5052),.B(g6210));
AND2X1 AND2_396 (.Y(g8699),.A(g7595),.B(g8579));
AND2X1 AND_tmp37 (.Y(ttmp37),.A(g1428),.B(g1432));
AND2X1 AND_tmp38 (.Y(ttmp38),.A(g1419),.B(ttmp37));
AND2X1 AND_tmp39 (.Y(I5689),.A(g1424),.B(ttmp38));
AND2X1 AND2_397 (.Y(g7820),.A(g1896),.B(g7479));
AND2X1 AND2_398 (.Y(g11021),.A(g448),.B(g10974));
AND2X1 AND2_399 (.Y(g5917),.A(g1044),.B(g5320));
AND2X1 AND2_400 (.Y(g6619),.A(g49),.B(g6156));
AND2X1 AND2_401 (.Y(g6318),.A(g1300),.B(g5949));
AND2X1 AND2_402 (.Y(g6872),.A(g1896),.B(g6389));
AND2X1 AND2_403 (.Y(g11320),.A(g11201),.B(g4379));
AND2X1 AND2_404 (.Y(g10514),.A(g10489),.B(g4580));
AND2X1 AND2_405 (.Y(g4006),.A(g201),.B(g3228));
AND2X1 AND2_406 (.Y(g9853),.A(g299),.B(g9771));
AND2X1 AND2_407 (.Y(g11274),.A(g4913),.B(g11197));
AND2X1 AND2_408 (.Y(g6193),.A(g2206),.B(g5151));
AND2X1 AND2_409 (.Y(g8119),.A(g6239),.B(g7890));
AND2X1 AND2_410 (.Y(g9420),.A(g1747),.B(g9030));
AND2X1 AND2_411 (.Y(g5233),.A(g1791),.B(g4492));
AND2X1 AND2_412 (.Y(g7581),.A(g7092),.B(g5420));
AND2X1 AND2_413 (.Y(g6549),.A(g5515),.B(g6175));
AND2X1 AND2_414 (.Y(g11464),.A(g11433),.B(g5446));
AND2X1 AND2_415 (.Y(g4801),.A(g516),.B(g3439));
AND2X1 AND2_416 (.Y(g6834),.A(g1365),.B(g6596));
AND2X1 AND2_417 (.Y(g4487),.A(g1718),.B(g3911));
AND2X1 AND2_418 (.Y(g2939),.A(g2411),.B(g1687));
AND2X1 AND2_419 (.Y(g7060),.A(g6739),.B(g5521));
AND2X1 AND2_420 (.Y(g5770),.A(g4466),.B(g5128));
AND2X1 AND2_421 (.Y(g5725),.A(g1580),.B(g5166));
AND2X1 AND2_422 (.Y(g11641),.A(g11615),.B(g7901));
AND2X1 AND2_423 (.Y(g2544),.A(g1341),.B(g1336));
AND2X1 AND2_424 (.Y(g11292),.A(g11252),.B(g4250));
AND2X1 AND2_425 (.Y(g5532),.A(g1681),.B(g4307));
AND2X1 AND2_426 (.Y(g11153),.A(g3771),.B(g10913));
AND2X1 AND2_427 (.Y(g9905),.A(g9872),.B(g9680));
AND2X1 AND2_428 (.Y(g7739),.A(g6957),.B(g3880));
AND2X1 AND2_429 (.Y(g6321),.A(g1284),.B(g5949));
AND2X1 AND2_430 (.Y(g8386),.A(g6085),.B(g8219));
AND2X1 AND_tmp40 (.Y(ttmp40),.A(g6764),.B(g8858));
AND2X1 AND_tmp41 (.Y(g8975),.A(g8089),.B(ttmp40));
AND2X1 AND2_431 (.Y(g2306),.A(g1223),.B(g1218));
AND2X1 AND2_432 (.Y(g6625),.A(g1218),.B(g6178));
AND2X1 AND2_433 (.Y(g7937),.A(g7606),.B(g4013));
AND2X1 AND2_434 (.Y(g10788),.A(g8303),.B(g10754));
AND2X1 AND2_435 (.Y(g10325),.A(g10248),.B(g3307));
AND2X1 AND2_436 (.Y(g8170),.A(g5270),.B(g7853));
AND2X1 AND2_437 (.Y(g5706),.A(g1574),.B(g5121));
AND2X1 AND2_438 (.Y(g2756),.A(g936),.B(g2081));
AND2X1 AND2_439 (.Y(g8821),.A(g8643),.B(g8751));
AND2X1 AND2_440 (.Y(g10946),.A(g5225),.B(g10827));
AND2X1 AND2_441 (.Y(g4169),.A(g2765),.B(g3066));
AND2X1 AND2_442 (.Y(g5029),.A(g1077),.B(g4521));
AND2X1 AND2_443 (.Y(g11164),.A(g4889),.B(g11112));
AND2X1 AND2_444 (.Y(g4007),.A(g2683),.B(g2276));
AND2X1 AND2_445 (.Y(g4059),.A(g1756),.B(g2796));
AND2X1 AND2_446 (.Y(g4868),.A(g1027),.B(g3914));
AND2X1 AND2_447 (.Y(g5675),.A(g131),.B(g5361));
AND2X1 AND2_448 (.Y(g4718),.A(g650),.B(g3343));
AND2X1 AND2_449 (.Y(g10682),.A(g10600),.B(g3863));
AND2X1 AND2_450 (.Y(g6687),.A(g5486),.B(g5840));
AND2X1 AND2_451 (.Y(g7704),.A(g682),.B(g7197));
AND2X1 AND2_452 (.Y(g4582),.A(g525),.B(g4055));
AND2X1 AND2_453 (.Y(g4261),.A(g1019),.B(g3914));
AND2X1 AND2_454 (.Y(g3422),.A(g225),.B(g3228));
AND2X1 AND2_455 (.Y(g5745),.A(g1549),.B(g5192));
AND2X1 AND2_456 (.Y(g8387),.A(g6086),.B(g8220));
AND2X1 AND2_457 (.Y(g7954),.A(g2874),.B(g7512));
AND2X1 AND2_458 (.Y(g11283),.A(g4966),.B(g11205));
AND2X1 AND2_459 (.Y(g8461),.A(g8298),.B(g7403));
AND2X1 AND2_460 (.Y(g10760),.A(g10695),.B(g10691));
AND2X1 AND2_461 (.Y(g11492),.A(g11480),.B(g4807));
AND2X1 AND_tmp42 (.Y(ttmp42),.A(g6626),.B(g5292));
AND2X1 AND_tmp43 (.Y(g7032),.A(g2965),.B(ttmp42));
AND2X1 AND2_462 (.Y(g8756),.A(g7431),.B(g8674));
AND2X1 AND2_463 (.Y(g9151),.A(g8967),.B(g6674));
AND2X1 AND2_464 (.Y(g6341),.A(g272),.B(g5885));
AND2X1 AND2_465 (.Y(g10506),.A(g10390),.B(g2135));
AND2X1 AND2_466 (.Y(g9648),.A(g16),.B(g9274));
AND2X1 AND2_467 (.Y(g7453),.A(g7148),.B(g2809));
AND2X1 AND2_468 (.Y(g6525),.A(g5995),.B(g3102));
AND2X1 AND2_469 (.Y(g6645),.A(g67),.B(g6202));
AND2X1 AND2_470 (.Y(g5707),.A(g1595),.B(g5122));
AND2X1 AND2_471 (.Y(g8046),.A(g7548),.B(g5128));
AND2X1 AND2_472 (.Y(g11091),.A(g833),.B(g10950));
AND2X1 AND2_473 (.Y(g11174),.A(g496),.B(g11112));
AND2X1 AND2_474 (.Y(g9010),.A(g6454),.B(g8930));
AND2X1 AND2_475 (.Y(g8403),.A(g6101),.B(g8239));
AND2X1 AND2_476 (.Y(g5201),.A(g1250),.B(g4721));
AND2X1 AND2_477 (.Y(g8841),.A(g8605),.B(g8704));
AND2X1 AND2_478 (.Y(g6879),.A(g1914),.B(g6407));
AND2X1 AND2_479 (.Y(g8763),.A(g7440),.B(g8680));
AND2X1 AND2_480 (.Y(g4502),.A(g2031),.B(g3938));
AND2X1 AND2_481 (.Y(g9839),.A(g9702),.B(g9742));
AND2X1 AND2_482 (.Y(g6358),.A(g5841),.B(g4441));
AND2X1 AND2_483 (.Y(g5575),.A(g1618),.B(g4501));
AND2X1 AND2_484 (.Y(g4940),.A(g3500),.B(g4440));
AND2X1 AND2_485 (.Y(g8107),.A(g6226),.B(g7882));
AND2X1 AND2_486 (.Y(g10240),.A(g10150),.B(g9103));
AND2X1 AND2_487 (.Y(g11192),.A(g5628),.B(g11066));
AND2X1 AND2_488 (.Y(g9618),.A(g910),.B(g9205));
AND2X1 AND2_489 (.Y(g5539),.A(g1684),.B(g4314));
AND2X1 AND2_490 (.Y(g8416),.A(g731),.B(g8151));
AND2X1 AND2_491 (.Y(g9693),.A(g275),.B(g9432));
AND2X1 AND2_492 (.Y(g11553),.A(g2683),.B(g11519));
AND2X1 AND2_493 (.Y(g8047),.A(g7557),.B(g5919));
AND2X1 AND2_494 (.Y(g5268),.A(g1098),.B(g4769));
AND2X1 AND2_495 (.Y(g9555),.A(g9107),.B(g3391));
AND2X1 AND2_496 (.Y(g6180),.A(g2190),.B(g5128));
AND2X1 AND2_497 (.Y(g6832),.A(g1383),.B(g6596));
AND2X1 AND2_498 (.Y(g10633),.A(g10600),.B(g3829));
AND2X1 AND2_499 (.Y(g7894),.A(g7617),.B(g3816));
AND2X1 AND2_500 (.Y(g8654),.A(g8529),.B(g4013));
AND2X1 AND2_501 (.Y(g9621),.A(g1179),.B(g9125));
AND2X1 AND2_502 (.Y(g6794),.A(g5819),.B(g4415));
AND2X1 AND2_503 (.Y(g9313),.A(g8876),.B(g5708));
AND2X1 AND2_504 (.Y(g4883),.A(g248),.B(g3946));
AND2X1 AND2_505 (.Y(g3412),.A(g219),.B(g3228));
AND2X1 AND2_506 (.Y(g7661),.A(g7127),.B(g2251));
AND2X1 AND_tmp44 (.Y(ttmp44),.A(g2369),.B(g591));
AND2X1 AND_tmp45 (.Y(g2800),.A(g2399),.B(ttmp44));
AND2X1 AND2_507 (.Y(g3389),.A(g207),.B(g3228));
AND2X1 AND2_508 (.Y(g3706),.A(g471),.B(g3268));
AND2X1 AND2_509 (.Y(g9908),.A(g9890),.B(g9782));
AND2X1 AND2_510 (.Y(g3429),.A(g231),.B(g3228));
AND2X1 AND2_511 (.Y(g6628),.A(g351),.B(g6182));
AND2X1 AND2_512 (.Y(g5470),.A(g1044),.B(g4222));
AND2X1 AND2_513 (.Y(g7526),.A(g7148),.B(g2868));
AND2X1 AND2_514 (.Y(g5897),.A(g2204),.B(g5354));
AND2X1 AND2_515 (.Y(g5025),.A(g1482),.B(g4640));
AND2X1 AND2_516 (.Y(g6204),.A(g3738),.B(g4921));
AND2X1 AND2_517 (.Y(g4048),.A(g1750),.B(g2790));
AND2X1 AND_tmp46 (.Y(ttmp46),.A(g6778),.B(g8849));
AND2X1 AND_tmp47 (.Y(g8935),.A(g8106),.B(ttmp46));
AND2X1 AND2_518 (.Y(g3281),.A(g766),.B(g2525));
AND2X1 AND2_519 (.Y(g9593),.A(g898),.B(g9205));
AND2X1 AND2_520 (.Y(g4827),.A(g213),.B(g3946));
AND2X1 AND2_521 (.Y(g10701),.A(g10620),.B(g10619));
AND2X1 AND2_522 (.Y(g10777),.A(g10733),.B(g3015));
AND2X1 AND2_523 (.Y(g8130),.A(g1936),.B(g7952));
AND2X1 AND2_524 (.Y(g9965),.A(g9955),.B(g9536));
AND2X1 AND2_525 (.Y(g3684),.A(g1710),.B(g3015));
AND2X1 AND2_526 (.Y(g11213),.A(g947),.B(g11157));
AND2X1 AND2_527 (.Y(g5006),.A(g1462),.B(g4640));
AND2X1 AND2_528 (.Y(g9933),.A(g9912),.B(g9624));
AND2X1 AND2_529 (.Y(g8554),.A(g8407),.B(g8020));
AND2X1 AND2_530 (.Y(g9641),.A(g913),.B(g9205));
AND2X1 AND2_531 (.Y(g6123),.A(g5630),.B(g4311));
AND2X1 AND2_532 (.Y(g6323),.A(g1235),.B(g5949));
AND2X1 AND2_533 (.Y(g10766),.A(g10646),.B(g4840));
AND2X1 AND2_534 (.Y(g6666),.A(g5301),.B(g5818));
AND2X1 AND2_535 (.Y(g4994),.A(g1504),.B(g4640));
AND2X1 AND2_536 (.Y(g5755),.A(g5103),.B(g5354));
AND2X1 AND2_537 (.Y(g11592),.A(g3717),.B(g11561));
AND2X1 AND2_538 (.Y(g6351),.A(g6210),.B(g5052));
AND2X1 AND2_539 (.Y(g6875),.A(g1905),.B(g6400));
AND2X1 AND2_540 (.Y(g4816),.A(g4070),.B(g2336));
AND2X1 AND2_541 (.Y(g9658),.A(g947),.B(g9240));
AND2X1 AND2_542 (.Y(g6530),.A(g6207),.B(g3829));
AND2X1 AND2_543 (.Y(g8366),.A(g8199),.B(g7265));
AND2X1 AND2_544 (.Y(g9835),.A(g9735),.B(g9785));
AND2X1 AND2_545 (.Y(g6655),.A(g5296),.B(g5812));
AND2X1 AND_tmp48 (.Y(ttmp48),.A(g3875),.B(g2733));
AND2X1 AND_tmp49 (.Y(g5445),.A(g4631),.B(ttmp48));
AND2X1 AND2_546 (.Y(g5173),.A(g3094),.B(g4676));
AND2X1 AND2_547 (.Y(g7970),.A(g7384),.B(g7703));
AND2X1 AND2_548 (.Y(g3098),.A(g2331),.B(g2198));
AND2X1 AND2_549 (.Y(g5491),.A(g1624),.B(g4262));
AND2X1 AND2_550 (.Y(g9271),.A(g6681),.B(g8949));
AND2X1 AND2_551 (.Y(g11152),.A(g369),.B(g10903));
AND2X1 AND2_552 (.Y(g9611),.A(g2651),.B(g9010));
AND2X1 AND2_553 (.Y(g6410),.A(g2804),.B(g5759));
AND2X1 AND2_554 (.Y(g10451),.A(g10444),.B(g3365));
AND2X1 AND2_555 (.Y(g4397),.A(g3475),.B(g2181));
AND2X1 AND2_556 (.Y(g7224),.A(g5398),.B(g6441));
AND2X1 AND2_557 (.Y(g5602),.A(g1624),.B(g4535));
AND2X1 AND2_558 (.Y(g4421),.A(g4112),.B(g2980));
AND2X1 AND2_559 (.Y(g6884),.A(g5569),.B(g6564));
AND2X1 AND2_560 (.Y(g6839),.A(g1397),.B(g6596));
AND2X1 AND2_561 (.Y(g8698),.A(g7591),.B(g8576));
AND2X1 AND_tmp50 (.Y(ttmp50),.A(g6368),.B(g8849));
AND2X1 AND_tmp51 (.Y(g8964),.A(g8255),.B(ttmp50));
AND2X1 AND2_562 (.Y(g8260),.A(g2775),.B(g7911));
AND2X1 AND2_563 (.Y(g11413),.A(g11354),.B(g10679));
AND2X1 AND2_564 (.Y(g4950),.A(g1415),.B(g4682));
AND2X1 AND2_565 (.Y(g5535),.A(g4327),.B(g3544));
AND2X1 AND2_566 (.Y(g7277),.A(g6772),.B(g731));
AND2X1 AND2_567 (.Y(g8463),.A(g8301),.B(g7410));
AND2X1 AND2_568 (.Y(g3268),.A(g466),.B(g2511));
AND2X1 AND2_569 (.Y(g10785),.A(g10728),.B(g5177));
AND2X1 AND2_570 (.Y(g6618),.A(g658),.B(g6016));
AND2X1 AND2_571 (.Y(g6235),.A(g569),.B(g5089));
AND2X1 AND2_572 (.Y(g10950),.A(g10788),.B(g6355));
AND2X1 AND2_573 (.Y(g4723),.A(g3626),.B(g2779));
AND2X1 AND2_574 (.Y(g8720),.A(g8601),.B(g7905));
AND2X1 AND2_575 (.Y(g6693),.A(g5494),.B(g5845));
AND2X1 AND2_576 (.Y(g11020),.A(g452),.B(g10974));
AND2X1 AND2_577 (.Y(g11583),.A(g1314),.B(g11541));
AND2X1 AND2_578 (.Y(g8118),.A(g1900),.B(g7941));
AND2X1 AND2_579 (.Y(g8167),.A(g5253),.B(g7853));
AND2X1 AND2_580 (.Y(g6334),.A(g1389),.B(g5904));
AND2X1 AND2_581 (.Y(g7892),.A(g7616),.B(g3815));
AND2X1 AND2_582 (.Y(g8652),.A(g8523),.B(g4013));
AND2X1 AND2_583 (.Y(g5721),.A(g1577),.B(g5143));
AND2X1 AND2_584 (.Y(g10367),.A(g10362),.B(g3375));
AND2X1 AND2_585 (.Y(g9901),.A(g9893),.B(g9392));
AND2X1 AND2_586 (.Y(g6792),.A(g290),.B(g5881));
AND2X1 AND2_587 (.Y(g11282),.A(g4958),.B(g11203));
AND2X1 AND2_588 (.Y(g7945),.A(g2847),.B(g7473));
AND2X1 AND_tmp52 (.Y(ttmp52),.A(g6764),.B(g8858));
AND2X1 AND_tmp53 (.Y(g8971),.A(g8081),.B(ttmp52));
AND2X1 AND2_589 (.Y(g11302),.A(g5508),.B(g11244));
AND2X1 AND2_590 (.Y(g4585),.A(g521),.B(g4060));
AND2X1 AND2_591 (.Y(g6621),.A(g52),.B(g6164));
AND2X1 AND2_592 (.Y(g5502),.A(g1932),.B(g4275));
AND2X1 AND2_593 (.Y(g11105),.A(g3634),.B(g10937));
AND2X1 AND2_594 (.Y(g7709),.A(g6856),.B(g4333));
AND2X1 AND2_595 (.Y(g8598),.A(g8471),.B(g7432));
AND2X1 AND2_596 (.Y(g7140),.A(g6069),.B(g6711));
AND2X1 AND2_597 (.Y(g9600),.A(g904),.B(g9205));
AND2X1 AND2_598 (.Y(g9864),.A(g1604),.B(g9778));
AND2X1 AND2_599 (.Y(g11640),.A(g11613),.B(g7900));
AND2X1 AND2_600 (.Y(g5188),.A(g4504),.B(g4496));
AND2X1 AND2_601 (.Y(g7435),.A(g7260),.B(g6572));
AND2X1 AND2_602 (.Y(g7876),.A(g7609),.B(g3790));
AND2X1 AND2_603 (.Y(g5030),.A(g1280),.B(g4523));
AND2X1 AND2_604 (.Y(g4058),.A(g2707),.B(g2276));
AND2X1 AND2_605 (.Y(g6776),.A(g5809),.B(g4390));
AND2X1 AND2_606 (.Y(g4890),.A(g630),.B(g4739));
AND2X1 AND2_607 (.Y(g2525),.A(g762),.B(g758));
AND2X1 AND2_608 (.Y(g10301),.A(g8892),.B(g10223));
AND2X1 AND2_609 (.Y(g4505),.A(g354),.B(g3586));
AND2X1 AND2_610 (.Y(g9623),.A(g17),.B(g9274));
AND2X1 AND2_611 (.Y(g10739),.A(g10676),.B(g3368));
AND2X1 AND2_612 (.Y(g11027),.A(g391),.B(g10974));
AND2X1 AND2_613 (.Y(g10738),.A(g10692),.B(g4840));
AND2X1 AND2_614 (.Y(g8687),.A(g8558),.B(g8036));
AND2X1 AND2_615 (.Y(g6360),.A(g302),.B(g5899));
AND2X1 AND2_616 (.Y(g9871),.A(g1564),.B(g9668));
AND2X1 AND2_617 (.Y(g5108),.A(g1801),.B(g4614));
AND2X1 AND2_618 (.Y(g11248),.A(g976),.B(g11071));
AND2X1 AND2_619 (.Y(g4992),.A(g1407),.B(g4682));
AND2X1 AND2_620 (.Y(g11552),.A(g2677),.B(g11519));
AND2X1 AND2_621 (.Y(g9651),.A(g944),.B(g9240));
AND2X1 AND2_622 (.Y(g11204),.A(g971),.B(g11083));
AND2X1 AND2_623 (.Y(g7824),.A(g1932),.B(g7479));
AND2X1 AND2_624 (.Y(g4480),.A(g1133),.B(g3905));
AND2X1 AND2_625 (.Y(g6179),.A(g5115),.B(g5354));
AND2X1 AND2_626 (.Y(g8710),.A(g7607),.B(g8595));
AND2X1 AND2_627 (.Y(g7590),.A(g7102),.B(g5425));
AND2X1 AND2_628 (.Y(g9384),.A(g968),.B(g9223));
AND2X1 AND2_629 (.Y(g3407),.A(g2561),.B(g3012));
AND2X1 AND2_630 (.Y(g9838),.A(g9700),.B(g9754));
AND2X1 AND2_631 (.Y(g3718),.A(g192),.B(g3164));
AND2X1 AND2_632 (.Y(g10661),.A(g10594),.B(g3015));
AND2X1 AND2_633 (.Y(g11380),.A(g11321),.B(g4285));
AND2X1 AND_tmp54 (.Y(ttmp54),.A(g6764),.B(g8858));
AND2X1 AND_tmp55 (.Y(g8879),.A(g8110),.B(ttmp54));
AND2X1 AND2_634 (.Y(g7930),.A(g7621),.B(g3110));
AND2X1 AND_tmp56 (.Y(ttmp56),.A(g6368),.B(g8828));
AND2X1 AND_tmp57 (.Y(g8962),.A(g8089),.B(ttmp56));
AND2X1 AND2_635 (.Y(g10715),.A(g2272),.B(g10630));
AND2X1 AND2_636 (.Y(g8659),.A(g8535),.B(g4013));
AND2X1 AND2_637 (.Y(g3015),.A(g2028),.B(g2191));
AND2X1 AND2_638 (.Y(g9643),.A(g950),.B(g9223));
AND2X1 AND2_639 (.Y(g9205),.A(g6454),.B(g8957));
AND2X1 AND2_640 (.Y(g5538),.A(g1669),.B(g4313));
AND2X1 AND2_641 (.Y(g4000),.A(g1744),.B(g2778));
AND2X1 AND2_642 (.Y(g4126),.A(g2701),.B(g3040));
AND2X1 AND2_643 (.Y(g4400),.A(g4088),.B(g3829));
AND2X1 AND2_644 (.Y(g2794),.A(I5886),.B(I5887));
AND2X1 AND2_645 (.Y(g4760),.A(g486),.B(g3393));
AND2X1 AND2_646 (.Y(g6238),.A(g572),.B(g5096));
AND2X1 AND2_647 (.Y(g10784),.A(g10727),.B(g5169));
AND2X1 AND2_648 (.Y(g8174),.A(g5284),.B(g7853));
AND2X1 AND2_649 (.Y(g6332),.A(g1374),.B(g5904));
AND2X1 AND2_650 (.Y(g5067),.A(g305),.B(g4811));
AND2X1 AND2_651 (.Y(g5418),.A(g1512),.B(g4344));
AND2X1 AND2_652 (.Y(g10297),.A(g8892),.B(g10211));
AND2X1 AND2_653 (.Y(g6353),.A(g299),.B(g5895));
AND2X1 AND2_654 (.Y(g11026),.A(g386),.B(g10974));
AND2X1 AND2_655 (.Y(g11212),.A(g944),.B(g11155));
NAND2X1 AND2_656 (.Y(g6744),.A(g4828),.B(g6151));
AND2X1 AND2_657 (.Y(g5493),.A(g1923),.B(g4265));
AND2X1 AND2_658 (.Y(g10671),.A(g10578),.B(g9431));
AND2X1 AND2_659 (.Y(g4383),.A(g2517),.B(g3829));
AND2X1 AND2_660 (.Y(g5256),.A(g4297),.B(g2779));
AND2X1 AND2_661 (.Y(g4220),.A(g105),.B(g3539));
AND2X1 AND2_662 (.Y(g8380),.A(g8252),.B(g4240));
AND2X1 AND2_663 (.Y(g7071),.A(g5916),.B(g6590));
AND2X1 AND2_664 (.Y(g4779),.A(g501),.B(g3427));
AND2X1 AND2_665 (.Y(g9613),.A(g1176),.B(g9125));
AND2X1 AND2_666 (.Y(g7705),.A(g6853),.B(g4328));
NAND2X1 AND2_667 (.Y(g9269),.A(g8933),.B(g3413));
AND2X1 AND2_668 (.Y(g5181),.A(g4520),.B(g4510));
AND2X1 AND2_669 (.Y(g4977),.A(g4567),.B(g4807));
AND2X1 AND2_670 (.Y(g7948),.A(g2855),.B(g7497));
AND2X1 AND2_671 (.Y(g11149),.A(g324),.B(g10930));
AND2X1 AND2_672 (.Y(g9862),.A(g1601),.B(g9777));
AND2X1 AND2_673 (.Y(g11387),.A(g11284),.B(g3629));
DFFX1 DFF_34 (.CK(CK1), .D(g8447), .Q(g1499));
DFFX1 DFF_35 (.CK(CK1), .D(g7789), .Q(g1044));
DFFX1 DFF_36 (.CK(CK1), .D(g8987), .Q(g1444));
DFFX1 DFF_37 (.CK(CK1), .D(g11179), .Q(g757));
DFFX1 DFF_38 (.CK(CK1), .D(g8436), .Q(g786));
DFFX1 DFF_39 (.CK(CK1), .D(g7344), .Q(g1543));
DFFX1 DFF_40 (.CK(CK1), .D(g11045), .Q(g552));
DFFX1 DFF_41 (.CK(CK1), .D(g5645), .Q(g315));
DFFX1 DFF_42 (.CK(CK1), .D(g7341), .Q(g1534));
DFFX1 DFF_43 (.CK(CK1), .D(g9338), .Q(g622));
DFFX1 DFF_44 (.CK(CK1), .D(g9354), .Q(g1927));
DFFX1 DFF_45 (.CK(CK1), .D(g11033), .Q(g1660));
DFFX1 DFF_46 (.CK(CK1), .D(g7765), .Q(g278));
DFFX1 DFF_47 (.CK(CK1), .D(g8989), .Q(g1436));
DFFX1 DFF_48 (.CK(CK1), .D(g8433), .Q(g718));
DFFX1 DFF_49 (.CK(CK1), .D(g7775), .Q(g76));
DFFX1 DFF_50 (.CK(CK1), .D(g11047), .Q(g554));
AND2X1 AND2_674 (.Y(g7955),.A(g2877),.B(g7516));
AND2X1 AND2_675 (.Y(g4161),.A(g2719),.B(g3060));
AND2X1 AND2_676 (.Y(g11148),.A(g2321),.B(g10913));
AND2X1 AND2_677 (.Y(g9712),.A(g1528),.B(g9490));
AND2X1 AND2_678 (.Y(g8931),.A(g8807),.B(g8164));
AND2X1 AND2_679 (.Y(g11097),.A(g378),.B(g10884));
AND2X1 AND_tmp58 (.Y(ttmp58),.A(g2733),.B(g3819));
AND2X1 AND_tmp59 (.Y(g5421),.A(g4631),.B(ttmp58));
AND2X1 AND2_680 (.Y(g11104),.A(g2963),.B(g10937));
AND2X1 AND2_681 (.Y(g5263),.A(g709),.B(g4761));
AND2X1 AND2_682 (.Y(g6092),.A(g1059),.B(g5320));
AND2X1 AND2_683 (.Y(g4999),.A(g1499),.B(g4640));
AND2X1 AND_tmp60 (.Y(ttmp60),.A(g2451),.B(g2446));
AND2X1 AND_tmp61 (.Y(ttmp61),.A(g2475),.B(ttmp60));
AND2X1 AND_tmp62 (.Y(I6338),.A(g2456),.B(ttmp61));
AND2X1 AND_tmp63 (.Y(ttmp63),.A(g632),.B(g6858));
AND2X1 AND_tmp64 (.Y(g7409),.A(g4976),.B(ttmp63));
AND2X1 AND2_684 (.Y(g4103),.A(g2683),.B(g2997));
AND2X1 AND_tmp65 (.Y(ttmp65),.A(g2456),.B(g2475));
AND2X1 AND_tmp66 (.Y(ttmp66),.A(g2446),.B(ttmp65));
AND2X1 AND_tmp67 (.Y(I6309),.A(g2451),.B(ttmp66));
AND2X1 AND2_685 (.Y(g6580),.A(g1801),.B(g5944));
AND2X1 AND2_686 (.Y(g5631),.A(g1056),.B(g4416));
AND2X1 AND2_687 (.Y(g9414),.A(g1730),.B(g9052));
NAND2X1 AND2_688 (.Y(g9660),.A(g1188),.B(g9125));
AND2X1 AND2_689 (.Y(g9946),.A(g9926),.B(g9392));
AND2X1 AND2_702 (.Y(g7822),.A(g1914),.B(g7479));
AND2X1 AND2_703 (.Y(g8123),.A(g1918),.B(g7946));
NAND2X1 AND2_704 (.Y(g11582),.A(g1311),.B(g11540));
AND2X1 AND2_705 (.Y(g4316),.A(g1965),.B(g3400));
AND2X1 AND2_706 (.Y(g10969),.A(g3625),.B(g10809));
AND2X1 AND2_707 (.Y(g5041),.A(g3983),.B(g4401));
AND2X1 AND2_708 (.Y(g9335),.A(g8975),.B(g5708));
AND2X1 AND2_709 (.Y(g9831),.A(g9727),.B(g9785));
AND2X1 AND2_710 (.Y(g4565),.A(g534),.B(g4010));
AND2X1 AND2_711 (.Y(g9422),.A(g1750),.B(g9030));
AND2X1 AND2_712 (.Y(g8648),.A(g4588),.B(g8511));
AND2X1 AND_tmp68 (.Y(ttmp68),.A(g6368),.B(g8858));
AND2X1 AND_tmp69 (.Y(g8875),.A(g8255),.B(ttmp68));
AND2X1 AND2_713 (.Y(g5168),.A(g1512),.B(g4679));
AND2X1 AND2_714 (.Y(g7895),.A(g7503),.B(g7036));
AND2X1 AND2_715 (.Y(g8655),.A(g8532),.B(g4013));
AND2X1 AND2_716 (.Y(g3396),.A(g213),.B(g3228));
AND2X1 AND2_717 (.Y(g4914),.A(g1062),.B(g4436));
AND2X1 AND2_718 (.Y(g9947),.A(g9927),.B(g9392));
AND2X1 AND2_719 (.Y(g5772),.A(g1555),.B(g5214));
AND2X1 AND2_720 (.Y(g6838),.A(g192),.B(g6596));
AND2X1 AND2_721 (.Y(g5531),.A(g1666),.B(g4306));
AND2X1 AND2_722 (.Y(g6795),.A(g5036),.B(g5878));
AND2X1 AND2_723 (.Y(g10503),.A(g10388),.B(g2135));
AND2X1 AND2_724 (.Y(g8010),.A(g7738),.B(g7413));
AND2X1 AND2_725 (.Y(g8410),.A(g713),.B(g8143));
AND2X1 AND2_726 (.Y(g6231),.A(g818),.B(g5608));
AND2X1 AND2_727 (.Y(g10581),.A(g10531),.B(g9453));
AND2X1 AND2_728 (.Y(g10450),.A(g10364),.B(g3359));
AND2X1 AND2_729 (.Y(g2804),.A(g2132),.B(g1891));
AND2X1 AND2_730 (.Y(g3418),.A(g2379),.B(g3012));
AND2X1 AND2_731 (.Y(g4820),.A(g186),.B(g3946));
AND2X1 AND2_732 (.Y(g9653),.A(g1185),.B(g9125));
AND2X1 AND2_733 (.Y(g6205),.A(g1515),.B(g5151));
AND2X1 AND2_734 (.Y(g10818),.A(g10730),.B(g4545));
AND2X1 AND2_735 (.Y(g8172),.A(g5275),.B(g7853));
AND2X1 AND2_736 (.Y(g10496),.A(g10429),.B(g3977));
AND2X1 AND2_737 (.Y(g5074),.A(g1771),.B(g4587));
AND2X1 AND2_738 (.Y(g9869),.A(g1558),.B(g9814));
AND2X1 AND2_739 (.Y(g9719),.A(g1543),.B(g9490));
AND2X1 AND2_740 (.Y(g10741),.A(g10635),.B(g4013));
AND2X1 AND2_741 (.Y(g3381),.A(g940),.B(g2756));
AND2X1 AND2_742 (.Y(g5863),.A(g5272),.B(g2173));
AND2X1 AND2_743 (.Y(g8693),.A(g3738),.B(g8509));
AND2X1 AND2_744 (.Y(g5480),.A(g4279),.B(g3519));
AND2X1 AND2_745 (.Y(g4581),.A(g3766),.B(g3254));
AND2X1 AND2_746 (.Y(g3685),.A(g1781),.B(g2981));
AND2X1 AND2_747 (.Y(g5569),.A(g4816),.B(g2338));
AND2X1 AND2_748 (.Y(g8555),.A(g8409),.B(g8025));
AND2X1 AND2_749 (.Y(g3263),.A(g2503),.B(g2328));
AND2X1 AND2_750 (.Y(g9364),.A(g965),.B(g9223));
AND2X1 AND2_751 (.Y(g4784),.A(g506),.B(g3432));
AND2X1 AND2_752 (.Y(g9454),.A(g8994),.B(g5708));
AND2X1 AND_tmp70 (.Y(ttmp70),.A(g2074),.B(g2077));
AND2X1 AND_tmp71 (.Y(ttmp71),.A(g2060),.B(ttmp70));
AND2X1 AND_tmp72 (.Y(I6331),.A(g2070),.B(ttmp71));
AND2X1 AND2_753 (.Y(g11299),.A(g5498),.B(g11243));
AND2X1 AND2_754 (.Y(g6983),.A(g6592),.B(g3105));
AND2X1 AND2_755 (.Y(g7958),.A(g736),.B(g7697));
AND2X1 AND2_756 (.Y(g4995),.A(g1474),.B(g4640));
AND2X1 AND2_757 (.Y(g4079),.A(g2765),.B(g2276));
AND2X1 AND2_758 (.Y(g2264),.A(g1771),.B(g1766));
AND2X1 AND2_759 (.Y(g2160),.A(g745),.B(g746));
AND2X1 AND2_760 (.Y(g3257),.A(g378),.B(g2496));
AND2X1 AND2_761 (.Y(g3101),.A(I6309),.B(I6310));
AND2X1 AND2_762 (.Y(g5000),.A(g1470),.B(g4640));
AND2X1 AND2_763 (.Y(g3301),.A(g1346),.B(g2544));
AND2X1 AND2_764 (.Y(g5126),.A(g3076),.B(g4638));
AND2X1 AND_tmp73 (.Y(ttmp73),.A(g1474),.B(g1478));
AND2X1 AND_tmp74 (.Y(ttmp74),.A(g1462),.B(ttmp73));
AND2X1 AND_tmp75 (.Y(I5084),.A(g1470),.B(ttmp74));
AND2X1 AND2_765 (.Y(g9412),.A(g1727),.B(g9052));
AND2X1 AND2_766 (.Y(g9389),.A(g1330),.B(g9151));
AND2X1 AND2_767 (.Y(g2379),.A(g744),.B(g743));
AND2X1 AND2_768 (.Y(g10706),.A(g10567),.B(g4840));
AND2X1 AND_tmp76 (.Y(ttmp76),.A(g10447),.B(g10446));
AND2X1 AND_tmp77 (.Y(I16145),.A(g10366),.B(ttmp76));
AND2X1 AND2_769 (.Y(g10597),.A(g10533),.B(g4359));
AND2X1 AND_tmp78 (.Y(ttmp78),.A(g6778),.B(g8849));
AND2X1 AND_tmp79 (.Y(g8965),.A(g8110),.B(ttmp78));
AND2X1 AND2_770 (.Y(g5608),.A(g814),.B(g4831));
AND2X1 AND2_771 (.Y(g5220),.A(g1083),.B(g4729));
AND2X1 AND2_772 (.Y(g10624),.A(g10545),.B(g4544));
AND2X1 AND2_773 (.Y(g10300),.A(g8892),.B(g10220));
AND2X1 AND2_774 (.Y(g5023),.A(g1071),.B(g4511));
AND2X1 AND2_775 (.Y(g4432),.A(g3723),.B(g1975));
AND2X1 AND2_776 (.Y(g4053),.A(g2701),.B(g2276));
AND2X1 AND2_777 (.Y(g8050),.A(g7596),.B(g5919));
AND2X1 AND2_778 (.Y(g5588),.A(g1639),.B(g4508));
AND2X1 AND_tmp80 (.Y(ttmp80),.A(g6074),.B(g2733));
AND2X1 AND_tmp81 (.Y(g6679),.A(g4631),.B(ttmp80));
AND2X1 AND2_779 (.Y(g9963),.A(g9953),.B(g9536));
AND2X1 AND2_780 (.Y(g3772),.A(g2542),.B(g3089));
AND2X1 AND2_781 (.Y(g5051),.A(g4432),.B(g2834));
AND2X1 AND2_782 (.Y(g6831),.A(g207),.B(g6596));
AND2X1 AND2_783 (.Y(g2981),.A(g1776),.B(g2264));
AND2X1 AND2_784 (.Y(g8724),.A(g8606),.B(g7910));
AND2X1 AND2_785 (.Y(g4157),.A(g2713),.B(g3055));
AND2X1 AND2_786 (.Y(g9707),.A(g1583),.B(g9474));
AND2X1 AND_tmp82 (.Y(ttmp82),.A(g6368),.B(g8858));
AND2X1 AND_tmp83 (.Y(g8878),.A(g8099),.B(ttmp82));
AND2X1 AND2_787 (.Y(g2132),.A(g1872),.B(g1882));
AND2X1 AND2_788 (.Y(g10763),.A(g10639),.B(g4840));
AND2X1 AND_tmp84 (.Y(ttmp84),.A(g8109),.B(g6475));
AND2X1 AND_tmp85 (.Y(g8289),.A(g6777),.B(ttmp84));
AND2X1 AND2_789 (.Y(g7898),.A(g7511),.B(g7041));
AND2X1 AND2_790 (.Y(g11271),.A(g5624),.B(g11191));
AND2X1 AND2_791 (.Y(g11461),.A(g11429),.B(g5446));
AND2X1 AND2_792 (.Y(g5732),.A(g1604),.B(g5176));
AND2X1 AND2_793 (.Y(g11145),.A(g315),.B(g10927));
AND2X1 AND2_794 (.Y(g11031),.A(g411),.B(g10974));
AND2X1 AND2_795 (.Y(g9865),.A(g1607),.B(g9780));
AND2X1 AND2_796 (.Y(g5944),.A(g1796),.B(g5233));
AND2X1 AND2_797 (.Y(g9715),.A(g1531),.B(g9490));
AND2X1 AND2_798 (.Y(g9604),.A(g1194),.B(g9111));
AND2X1 AND2_799 (.Y(g8799),.A(g8647),.B(g8727));
AND2X1 AND2_800 (.Y(g11198),.A(g4919),.B(g11069));
AND2X1 AND2_801 (.Y(g6873),.A(g3263),.B(g6557));
AND2X1 AND2_802 (.Y(g6632),.A(g61),.B(g6190));
AND2X1 AND2_803 (.Y(g6095),.A(g1062),.B(g5320));
AND2X1 AND2_804 (.Y(g3863),.A(g3323),.B(g2728));
AND2X1 AND2_805 (.Y(g9833),.A(g9729),.B(g9785));
AND2X1 AND2_806 (.Y(g6653),.A(g70),.B(g6213));
AND2X1 AND2_807 (.Y(g6102),.A(g1038),.B(g5320));
AND2X1 AND2_808 (.Y(g7819),.A(g1887),.B(g7479));
AND2X1 AND2_809 (.Y(g11393),.A(g11280),.B(g7916));
AND2X1 AND2_810 (.Y(g2511),.A(g461),.B(g456));
AND2X1 AND2_811 (.Y(g7088),.A(g2331),.B(g6737));
AND2X1 AND2_812 (.Y(g9584),.A(g2726),.B(g9173));
AND2X1 AND2_813 (.Y(g9896),.A(g9883),.B(g9624));
AND2X1 AND_tmp86 (.Y(ttmp86),.A(g3792),.B(g7980));
AND2X1 AND_tmp87 (.Y(g8209),.A(g4094),.B(ttmp86));
AND2X1 AND2_814 (.Y(g6752),.A(g6187),.B(g2343));
AND2X1 AND2_815 (.Y(g4778),.A(g421),.B(g3426));
AND2X1 AND2_816 (.Y(g11161),.A(g1969),.B(g10937));
AND2X1 AND2_817 (.Y(g9268),.A(g6681),.B(g8947));
AND2X1 AND2_818 (.Y(g5681),.A(g135),.B(g5361));
AND2X1 AND2_819 (.Y(g7951),.A(g2868),.B(g7505));
AND2X1 AND2_820 (.Y(g9419),.A(g1744),.B(g9030));
AND2X1 AND2_821 (.Y(g10268),.A(g10183),.B(g3307));
AND2X1 AND2_822 (.Y(g5533),.A(g1724),.B(g4308));
AND2X1 AND2_823 (.Y(g9052),.A(g8936),.B(g7192));
AND2X1 AND2_824 (.Y(g6786),.A(g178),.B(g5919));
AND2X1 AND2_825 (.Y(g10670),.A(g10571),.B(g9091));
AND2X1 AND2_826 (.Y(g11087),.A(g829),.B(g10950));
AND2X1 AND2_827 (.Y(g4949),.A(g3505),.B(g4449));
AND2X1 AND2_828 (.Y(g6364),.A(g5851),.B(g4454));
AND2X1 AND2_829 (.Y(g7825),.A(g1941),.B(g7479));
AND2X1 AND2_830 (.Y(g3400),.A(g115),.B(g3164));
AND2X1 AND2_831 (.Y(g4998),.A(g1304),.B(g4485));
AND2X1 AND2_832 (.Y(g10667),.A(g10576),.B(g9427));
AND2X1 AND2_833 (.Y(g7136),.A(g6050),.B(g6704));
AND2X1 AND2_834 (.Y(g6532),.A(g339),.B(g6057));
AND2X1 AND2_835 (.Y(g9385),.A(g1324),.B(g9151));
AND2X1 AND_tmp88 (.Y(ttmp88),.A(g1444),.B(g1448));
AND2X1 AND_tmp89 (.Y(ttmp89),.A(g1436),.B(ttmp88));
AND2X1 AND_tmp90 (.Y(I5690),.A(g1440),.B(ttmp89));
AND2X1 AND2_836 (.Y(g4484),.A(g1137),.B(g3909));
AND2X1 AND2_837 (.Y(g9897),.A(g9884),.B(g9624));
AND2X1 AND2_838 (.Y(g9425),.A(g1753),.B(g9030));
AND2X1 AND2_839 (.Y(g3383),.A(g186),.B(g3228));
AND2X1 AND2_840 (.Y(g5601),.A(g1035),.B(g4375));
AND2X1 AND2_841 (.Y(g7943),.A(g2840),.B(g7467));
AND2X1 AND2_842 (.Y(g11171),.A(g481),.B(g11112));
AND2X1 AND2_843 (.Y(g3423),.A(I6630),.B(I6631));
AND2X1 AND2_844 (.Y(g7230),.A(g6064),.B(g6444));
AND2X1 AND2_845 (.Y(g4952),.A(g1648),.B(g4457));
AND2X1 AND2_846 (.Y(g8736),.A(g7439),.B(g8635));
AND2X1 AND2_847 (.Y(g6787),.A(g266),.B(g5875));
AND2X1 AND_tmp91 (.Y(ttmp91),.A(g6778),.B(g8849));
AND2X1 AND_tmp92 (.Y(g8968),.A(g8089),.B(ttmp91));
AND2X1 AND2_848 (.Y(g10306),.A(g10214),.B(g9082));
AND2X1 AND2_849 (.Y(g9331),.A(g8972),.B(g5708));
AND2X1 AND2_850 (.Y(g11459),.A(g11427),.B(g5446));
AND2X1 AND2_851 (.Y(g4561),.A(g538),.B(g4003));
AND2X1 AND2_852 (.Y(g11425),.A(g11350),.B(g10899));
AND2X1 AND2_853 (.Y(g11458),.A(g11426),.B(g5446));
AND2X1 AND2_854 (.Y(g5739),.A(g1607),.B(g5185));
AND2X1 AND2_855 (.Y(g7496),.A(g7148),.B(g2840));
AND2X1 AND2_856 (.Y(g4986),.A(g1411),.B(g4682));
AND2X1 AND2_857 (.Y(g11010),.A(g5187),.B(g10827));
AND2X1 AND2_858 (.Y(g3999),.A(g1741),.B(g2777));
AND2X1 AND2_859 (.Y(g8175),.A(g5291),.B(g7853));
AND2X1 AND2_860 (.Y(g8722),.A(g8604),.B(g7908));
AND2X1 AND2_861 (.Y(g4764),.A(g411),.B(g3404));
AND2X1 AND2_862 (.Y(g7137),.A(g5590),.B(g6361));
AND2X1 AND2_863 (.Y(g7891),.A(g7471),.B(g7028));
AND2X1 AND2_864 (.Y(g8651),.A(g8520),.B(g4013));
AND2X1 AND2_865 (.Y(g5479),.A(g1845),.B(g4243));
AND2X1 AND2_866 (.Y(g11599),.A(g1341),.B(g11572));
AND2X1 AND2_867 (.Y(g6684),.A(g5314),.B(g5836));
AND2X1 AND2_868 (.Y(g6745),.A(g5605),.B(g6158));
AND2X1 AND2_869 (.Y(g6639),.A(g357),.B(g6196));
AND2X1 AND2_870 (.Y(g10937),.A(g4822),.B(g10822));
AND2X1 AND2_871 (.Y(g3696),.A(g1713),.B(g3015));
AND2X1 AND2_872 (.Y(g4503),.A(g654),.B(g3943));
AND2X1 AND2_873 (.Y(g6791),.A(g269),.B(g5880));
AND2X1 AND2_874 (.Y(g5190),.A(g1245),.B(g4716));
AND2X1 AND2_875 (.Y(g5390),.A(g3220),.B(g4819));
AND2X1 AND2_876 (.Y(g8384),.A(g8180),.B(g3397));
AND2X1 AND2_877 (.Y(g4224),.A(g1092),.B(g3638));
AND2X1 AND2_878 (.Y(g5501),.A(g1672),.B(g4273));
AND2X1 AND2_879 (.Y(g9173),.A(g8968),.B(g6674));
AND2X1 AND2_880 (.Y(g6759),.A(g148),.B(g5919));
AND2X1 AND2_881 (.Y(g8838),.A(g8602),.B(g8702));
AND2X1 AND2_882 (.Y(g8024),.A(g7394),.B(g4337));
AND2X1 AND2_883 (.Y(g10666),.A(g10575),.B(g9424));
AND2X1 AND2_884 (.Y(g11158),.A(g309),.B(g10935));
AND2X1 AND2_885 (.Y(g9602),.A(g2650),.B(g9010));
AND2X1 AND2_886 (.Y(g5704),.A(g143),.B(g5361));
AND2X1 AND2_887 (.Y(g4617),.A(g3275),.B(g3879));
AND2X1 AND2_888 (.Y(g11561),.A(g11518),.B(g3015));
AND2X1 AND2_889 (.Y(g9868),.A(g1555),.B(g9812));
AND2X1 AND2_890 (.Y(g11295),.A(g5475),.B(g11239));
AND2X1 AND2_891 (.Y(g11144),.A(g305),.B(g10926));
AND2X1 AND2_892 (.Y(g9718),.A(g1540),.B(g9490));
AND2X1 AND2_893 (.Y(g3434),.A(g237),.B(g3228));
AND2X1 AND2_894 (.Y(g4987),.A(g1440),.B(g4682));
AND2X1 AND2_895 (.Y(g4771),.A(g496),.B(g3416));
AND2X1 AND2_896 (.Y(g5250),.A(g1270),.B(g4748));
AND2X1 AND2_897 (.Y(g6098),.A(g1065),.B(g5320));
AND2X1 AND2_898 (.Y(g9582),.A(g2725),.B(g9173));
NAND2X1 AND2_899 (.Y(g6833),.A(g186),.B(g6596));
AND2X1 AND2_900 (.Y(g3533),.A(g1981),.B(g2892));
AND2X1 AND2_901 (.Y(g4892),.A(g632),.B(g4739));
AND2X1 AND2_902 (.Y(g8104),.A(g6218),.B(g7880));
AND2X1 AND2_903 (.Y(g9415),.A(g1733),.B(g9052));
NAND2X1 AND2_904 (.Y(g8499),.A(g8377),.B(g4737));
AND2X1 AND2_905 (.Y(g9664),.A(g1191),.B(g9125));
AND2X1 AND2_906 (.Y(g10740),.A(g10676),.B(g3384));
AND2X1 AND2_907 (.Y(g2534),.A(g798),.B(g794));
AND2X1 AND2_908 (.Y(g8754),.A(g7420),.B(g8667));
AND2X1 AND2_909 (.Y(g9721),.A(g9413),.B(g4785));
NAND2X1 AND2_910 (.Y(g6162),.A(g3584),.B(g5200));
AND2X1 AND2_911 (.Y(g4991),.A(g1508),.B(g4640));
AND2X1 AND2_912 (.Y(g6362),.A(g5846),.B(g4450));
AND2X1 AND_tmp93 (.Y(ttmp93),.A(g2719),.B(g2765));
AND2X1 AND_tmp94 (.Y(ttmp94),.A(g2707),.B(ttmp93));
AND2X1 AND_tmp95 (.Y(I6631),.A(g2713),.B(ttmp94));
AND2X1 AND2_913 (.Y(g10685),.A(g10608),.B(g3863));
AND2X1 AND2_914 (.Y(g4340),.A(g1153),.B(g3715));
AND2X1 AND2_915 (.Y(g11023),.A(g440),.B(g10974));
AND2X1 AND2_916 (.Y(g8044),.A(g7598),.B(g5919));
AND2X1 AND2_917 (.Y(g11224),.A(g968),.B(g11056));
AND2X1 AND2_918 (.Y(g11571),.A(g2018),.B(g11561));
AND2X1 AND2_919 (.Y(g4959),.A(g1520),.B(g4682));
AND2X1 AND2_920 (.Y(g10334),.A(g10265),.B(g3307));
AND2X1 AND2_921 (.Y(g5626),.A(g1633),.B(g4557));
AND2X1 AND2_922 (.Y(g9940),.A(g9920),.B(g9367));
AND2X1 AND2_923 (.Y(g4876),.A(g1086),.B(g3638));
AND2X1 AND2_924 (.Y(g6728),.A(g6250),.B(g4318));
AND2X1 AND2_925 (.Y(g6730),.A(g1872),.B(g6128));
AND2X1 AND2_926 (.Y(g9689),.A(g263),.B(g9432));
AND2X1 AND2_927 (.Y(g10762),.A(g10635),.B(g4840));
AND2X1 AND2_928 (.Y(g6070),.A(g1050),.B(g5320));
AND2X1 AND2_929 (.Y(g9428),.A(g1756),.B(g9030));
AND2X1 AND2_930 (.Y(g9030),.A(g8935),.B(g7192));
AND2X1 AND2_931 (.Y(g9430),.A(g1759),.B(g9030));
AND2X1 AND2_932 (.Y(g8927),.A(g7872),.B(g8807));
AND2X1 AND2_933 (.Y(g7068),.A(g5912),.B(g6586));
AND2X1 AND2_934 (.Y(g8014),.A(g7740),.B(g7419));
AND2X1 AND2_935 (.Y(g11392),.A(g11278),.B(g7914));
AND2X1 AND2_936 (.Y(g5782),.A(g1558),.B(g5223));
AND2X1 AND2_937 (.Y(g9910),.A(g9892),.B(g9809));
AND2X1 AND2_938 (.Y(g4824),.A(g774),.B(g4099));
AND2X1 AND2_939 (.Y(g6331),.A(g201),.B(g5904));
AND2X1 AND2_940 (.Y(g4236),.A(g1098),.B(g3638));
AND2X1 AND2_941 (.Y(g11559),.A(g2719),.B(g11519));
AND2X1 AND2_942 (.Y(g9609),.A(g907),.B(g9205));
AND2X1 AND2_943 (.Y(g11558),.A(g2713),.B(g11519));
AND2X1 AND2_944 (.Y(g6087),.A(g1056),.B(g5320));
AND2X1 AND2_945 (.Y(g4877),.A(g243),.B(g3946));
AND2X1 AND2_946 (.Y(g5526),.A(g1950),.B(g4294));
AND2X1 AND2_947 (.Y(g10751),.A(g10646),.B(g4013));
AND2X1 AND2_948 (.Y(g10772),.A(g10655),.B(g4840));
AND2X1 AND2_949 (.Y(g8135),.A(g1945),.B(g7956));
AND2X1 AND2_950 (.Y(g11544),.A(g11515),.B(g10584));
AND2X1 AND2_951 (.Y(g5084),.A(g1776),.B(g4591));
AND2X1 AND2_952 (.Y(g8382),.A(g6077),.B(g8213));
AND2X1 AND2_953 (.Y(g10230),.A(g8892),.B(g10145));
AND2X1 AND2_954 (.Y(g5484),.A(g1896),.B(g4256));
AND2X1 AND2_955 (.Y(g7241),.A(g6772),.B(g6172));
AND2X1 AND2_956 (.Y(g3942),.A(g219),.B(g3164));
AND2X1 AND2_957 (.Y(g10638),.A(g10608),.B(g3829));
AND2X1 AND2_958 (.Y(g4064),.A(g1759),.B(g2799));
AND2X1 AND2_959 (.Y(g9365),.A(g1321),.B(g9151));
AND2X1 AND2_960 (.Y(g9861),.A(g9738),.B(g9579));
AND2X1 AND2_961 (.Y(g8749),.A(g7604),.B(g8660));
AND2X1 AND2_962 (.Y(g11255),.A(g456),.B(g11075));
AND2X1 AND2_963 (.Y(g11189),.A(g5616),.B(g11064));
AND2X1 AND2_964 (.Y(g10510),.A(g10393),.B(g2135));
AND2X1 AND_tmp96 (.Y(ttmp96),.A(g6368),.B(g8828));
AND2X1 AND_tmp97 (.Y(g8947),.A(g8056),.B(ttmp96));
AND2X1 AND2_965 (.Y(g2917),.A(g2424),.B(g1657));
AND2X1 AND2_966 (.Y(g5919),.A(g5216),.B(g2965));
AND2X1 AND2_967 (.Y(g11188),.A(g5604),.B(g11063));
AND2X1 AND2_968 (.Y(g9846),.A(g287),.B(g9764));
AND2X1 AND2_969 (.Y(g7818),.A(g1878),.B(g7479));
AND2X1 AND2_970 (.Y(g11460),.A(g11428),.B(g5446));
AND2X1 AND2_971 (.Y(g5276),.A(g736),.B(g4780));
AND2X1 AND2_972 (.Y(g11030),.A(g406),.B(g10974));
AND2X1 AND2_973 (.Y(g11093),.A(g841),.B(g10950));
AND2X1 AND2_974 (.Y(g7893),.A(g7478),.B(g7031));
AND2X1 AND2_975 (.Y(g8653),.A(g8526),.B(g4013));
AND2X1 AND2_976 (.Y(g10442),.A(g10311),.B(g2135));
AND2X1 AND2_977 (.Y(g6535),.A(g345),.B(g6063));
AND2X1 AND2_978 (.Y(g8102),.A(g6209),.B(g7878));
AND2X1 AND_tmp98 (.Y(ttmp98),.A(g1504),.B(g1508));
AND2X1 AND_tmp99 (.Y(ttmp99),.A(g1490),.B(ttmp98));
AND2X1 AND_tmp100 (.Y(I5085),.A(g1494),.B(ttmp99));
AND2X1 AND2_979 (.Y(g5004),.A(g1296),.B(g4499));
AND2X1 AND2_980 (.Y(g3912),.A(g207),.B(g3164));
AND2X1 AND2_981 (.Y(g7186),.A(g2503),.B(g6403));
AND2X1 AND2_982 (.Y(g4489),.A(g348),.B(g3586));
AND2X1 AND2_983 (.Y(g9662),.A(g2094),.B(g9292));
AND2X1 AND2_984 (.Y(g9418),.A(g1741),.B(g9052));
AND2X1 AND2_985 (.Y(g11218),.A(g959),.B(g11053));
AND2X1 AND2_986 (.Y(g4471),.A(g1121),.B(g3862));
AND2X1 AND2_987 (.Y(g10746),.A(g10643),.B(g4013));
AND2X1 AND2_988 (.Y(g7125),.A(g1212),.B(g6648));
AND2X1 AND2_989 (.Y(g7821),.A(g1905),.B(g7479));
AND2X1 AND2_990 (.Y(g6246),.A(g178),.B(g5361));
AND2X1 AND2_991 (.Y(g9256),.A(g6689),.B(g8963));
AND2X1 AND2_992 (.Y(g8042),.A(g7533),.B(g5128));
AND2X1 AND2_993 (.Y(g10237),.A(g10145),.B(g9100));
AND2X1 AND2_994 (.Y(g7939),.A(g2829),.B(g7460));
AND2X1 AND2_995 (.Y(g8786),.A(g8638),.B(g8716));
AND2X1 AND2_996 (.Y(g10684),.A(g10604),.B(g3863));
AND2X1 AND2_997 (.Y(g11455),.A(g11435),.B(g5446));
AND2X1 AND2_998 (.Y(g8364),.A(g658),.B(g8235));
AND2X1 AND_tmp101 (.Y(ttmp101),.A(g2557),.B(g1814));
AND2X1 AND_tmp102 (.Y(g2990),.A(g2061),.B(ttmp101));
AND2X1 AND2_999 (.Y(g9847),.A(g290),.B(g9766));
AND2X1 AND2_1000 (.Y(g8054),.A(g7584),.B(g5919));
AND2X1 AND2_1001 (.Y(g5617),.A(g1050),.B(g4391));
AND2X1 AND2_1002 (.Y(g6502),.A(g5981),.B(g3095));
AND2X1 AND2_1003 (.Y(g5789),.A(g1561),.B(g5232));
AND2X1 AND2_1004 (.Y(g4009),.A(g1747),.B(g2789));
AND2X1 AND2_1005 (.Y(g11277),.A(g4920),.B(g11199));
AND2X1 AND2_1006 (.Y(g6940),.A(g6472),.B(g1945));
AND2X1 AND2_1007 (.Y(g7061),.A(g790),.B(g6760));
AND2X1 AND2_1008 (.Y(g11595),.A(g1336),.B(g11575));
AND2X1 AND2_1009 (.Y(g5771),.A(g1534),.B(g5213));
AND2X1 AND2_1010 (.Y(g8553),.A(g8405),.B(g8015));
AND2X1 AND2_1011 (.Y(g4836),.A(g643),.B(g3520));
AND2X1 AND2_1012 (.Y(g5547),.A(g1733),.B(g4326));
AND2X1 AND2_1013 (.Y(g6216),.A(g2232),.B(g5151));
AND2X1 AND2_1014 (.Y(g4967),.A(g1515),.B(g4682));
AND2X1 AND2_1015 (.Y(g6671),.A(g342),.B(g6227));
AND2X1 AND2_1016 (.Y(g7200),.A(g3098),.B(g6418));
AND2X1 AND2_1017 (.Y(g3661),.A(g382),.B(g3257));
AND2X1 AND2_1018 (.Y(g7046),.A(g5892),.B(g6570));
AND2X1 AND2_1019 (.Y(g4229),.A(g999),.B(g3914));
AND2X1 AND2_1020 (.Y(g8389),.A(g6091),.B(g8225));
AND2X1 AND2_1021 (.Y(g6430),.A(g5044),.B(g5791));
AND2X1 AND2_1022 (.Y(g8706),.A(g7602),.B(g8589));
AND2X1 AND2_1023 (.Y(g4993),.A(g1448),.B(g4682));
AND2X1 AND2_1024 (.Y(g6247),.A(g127),.B(g5361));
AND2X1 AND2_1025 (.Y(g9257),.A(g6689),.B(g8964));
AND2X1 AND2_1026 (.Y(g11170),.A(g525),.B(g11112));
AND2X1 AND2_1027 (.Y(g7145),.A(g6082),.B(g6718));
AND2X1 AND2_1028 (.Y(g5738),.A(g1586),.B(g5184));
AND2X1 AND2_1029 (.Y(g6826),.A(g225),.B(g6596));
AND2X1 AND2_1030 (.Y(g7191),.A(g6343),.B(g4323));
AND2X1 AND2_1031 (.Y(g3998),.A(g2677),.B(g2276));
AND2X1 AND2_1032 (.Y(g6741),.A(g3284),.B(g6141));
AND2X1 AND2_1033 (.Y(g5478),.A(g1905),.B(g4242));
AND2X1 AND2_1034 (.Y(g11167),.A(g538),.B(g11112));
AND2X1 AND2_1035 (.Y(g11194),.A(g5637),.B(g11067));
AND2X1 AND2_1036 (.Y(g11589),.A(g1333),.B(g11548));
AND2X1 AND2_1037 (.Y(g6638),.A(g64),.B(g6195));
AND2X1 AND2_1038 (.Y(g4921),.A(g2779),.B(g4431));
AND2X1 AND2_1039 (.Y(g7536),.A(g7148),.B(g2877));
AND2X1 AND2_1040 (.Y(g9585),.A(g889),.B(g8995));
AND2X1 AND2_1041 (.Y(g2957),.A(g2424),.B(g1663));
AND2X1 AND2_1042 (.Y(g11588),.A(g1330),.B(g11547));
AND2X1 AND2_1043 (.Y(g5690),.A(g1567),.B(g5112));
AND2X1 AND2_1044 (.Y(g6883),.A(g1923),.B(g6413));
AND2X1 AND2_1045 (.Y(g4837),.A(g1068),.B(g3638));
AND2X1 AND_tmp103 (.Y(ttmp103),.A(g6368),.B(g8849));
AND2X1 AND_tmp104 (.Y(g8963),.A(g8056),.B(ttmp103));
AND2X1 AND2_1046 (.Y(g8791),.A(g8641),.B(g8721));
AND2X1 AND2_1047 (.Y(g6217),.A(g563),.B(g5073));
AND2X1 AND_tmp105 (.Y(ttmp105),.A(g2381),.B(g2395));
AND2X1 AND_tmp106 (.Y(ttmp106),.A(g2082),.B(ttmp105));
AND2X1 AND_tmp107 (.Y(I6316),.A(g2087),.B(ttmp106));
AND2X1 AND2_1048 (.Y(g11022),.A(g444),.B(g10974));
AND2X1 AND2_1049 (.Y(g5915),.A(g4168),.B(g4977));
AND2X1 AND2_1050 (.Y(g4788),.A(g511),.B(g3436));
AND2X1 AND2_1051 (.Y(g8759),.A(g7437),.B(g8677));
AND2X1 AND2_1052 (.Y(g5110),.A(g1806),.B(g4618));
AND2X1 AND2_1053 (.Y(g11254),.A(g986),.B(g11073));
AND2X1 AND2_1054 (.Y(g6827),.A(g219),.B(g6596));
AND2X1 AND_tmp108 (.Y(ttmp108),.A(g6368),.B(g8828));
AND2X1 AND_tmp109 (.Y(g8957),.A(g8081),.B(ttmp108));
AND2X1 AND2_1055 (.Y(g6333),.A(g197),.B(g5904));
AND2X1 AND2_1056 (.Y(g8049),.A(g7567),.B(g5919));
AND2X1 AND2_1057 (.Y(g4392),.A(g3273),.B(g3829));
AND2X1 AND2_1058 (.Y(g9856),.A(g1592),.B(g9773));
AND2X1 AND2_1059 (.Y(g9411),.A(g1724),.B(g9052));
AND2X1 AND2_1060 (.Y(g5002),.A(g1494),.B(g4640));
AND2X1 AND2_1061 (.Y(g11101),.A(g857),.B(g10950));
AND2X1 AND2_1062 (.Y(g11177),.A(g511),.B(g11112));
AND2X1 AND2_1063 (.Y(g11560),.A(g2765),.B(g11519));
AND2X1 AND2_1064 (.Y(g8098),.A(g6201),.B(g7852));
AND2X1 AND2_1065 (.Y(g3970),.A(g225),.B(g3164));
AND2X1 AND2_1066 (.Y(g4941),.A(g1038),.B(g4451));
AND2X1 AND2_1067 (.Y(g10453),.A(g10437),.B(g3395));
AND2X1 AND2_1068 (.Y(g5877),.A(g4921),.B(g639));
AND2X1 AND2_1069 (.Y(g6662),.A(g366),.B(g6220));
AND2X1 AND2_1070 (.Y(g7935),.A(g2821),.B(g7454));
AND2X1 AND2_1071 (.Y(g6067),.A(g1047),.B(g5320));
AND2X1 AND_tmp110 (.Y(ttmp110),.A(g2434),.B(g2438));
AND2X1 AND_tmp111 (.Y(ttmp111),.A(g2406),.B(ttmp110));
AND2X1 AND_tmp112 (.Y(I6317),.A(g2420),.B(ttmp111));
AND2X1 AND2_1072 (.Y(g9863),.A(g9740),.B(g9576));
AND2X1 AND_tmp113 (.Y(ttmp113),.A(g2249),.B(g2254));
AND2X1 AND_tmp114 (.Y(ttmp114),.A(g174),.B(ttmp113));
AND2X1 AND_tmp115 (.Y(I5886),.A(g170),.B(ttmp114));
AND2X1 AND2_1073 (.Y(g6994),.A(g6758),.B(g3829));
AND2X1 AND2_1074 (.Y(g9713),.A(g1589),.B(g9474));
AND2X1 AND2_1075 (.Y(g4431),.A(g2268),.B(g3533));
AND2X1 AND2_1076 (.Y(g4252),.A(g1007),.B(g3914));
AND2X1 AND2_1077 (.Y(g11166),.A(g542),.B(g11112));
AND2X1 AND2_1078 (.Y(g7130),.A(g6041),.B(g6697));
AND2X1 AND2_1079 (.Y(g11009),.A(g5179),.B(g10827));
AND2X1 AND2_1080 (.Y(g7542),.A(g7148),.B(g2885));
AND2X1 AND2_1081 (.Y(g8019),.A(g7386),.B(g4332));
AND2X1 AND2_1082 (.Y(g11008),.A(g5171),.B(g10827));
AND2X1 AND2_1083 (.Y(g3516),.A(g1209),.B(g3015));
AND2X1 AND2_1084 (.Y(g8052),.A(g7573),.B(g5128));
AND2X1 AND2_1085 (.Y(g3987),.A(g243),.B(g3164));
AND2X1 AND2_1086 (.Y(g4765),.A(g491),.B(g3405));
AND2X1 AND2_1087 (.Y(g11555),.A(g2695),.B(g11519));
AND2X1 AND2_1088 (.Y(g9857),.A(g9734),.B(g9569));
AND2X1 AND2_1089 (.Y(g8728),.A(g8610),.B(g7915));
AND2X1 AND2_1090 (.Y(g8730),.A(g8613),.B(g7917));
AND2X1 AND2_1091 (.Y(g8185),.A(g664),.B(g7997));
AND2X1 AND2_1092 (.Y(g5194),.A(g1610),.B(g4717));
AND2X1 AND2_1093 (.Y(g8385),.A(g6084),.B(g8218));
AND2X1 AND2_1094 (.Y(g4610),.A(g3804),.B(g2212));
AND2X1 AND2_1095 (.Y(g7902),.A(g7661),.B(g6587));
AND2X1 AND2_1096 (.Y(g4073),.A(g3200),.B(g3222));
AND2X1 AND2_1097 (.Y(g8070),.A(g682),.B(g7826));
AND2X1 AND2_1098 (.Y(g5731),.A(g1583),.B(g5175));
AND2X1 AND2_1099 (.Y(g11238),.A(g5474),.B(g11110));
AND2X1 AND2_1100 (.Y(g4473),.A(g1125),.B(g3874));
AND2X1 AND2_1101 (.Y(g8470),.A(g8308),.B(g7427));
AND2X1 AND2_1102 (.Y(g5489),.A(g4287),.B(g3521));
AND2X1 AND2_1103 (.Y(g3991),.A(g1738),.B(g2774));
AND2X1 AND_tmp116 (.Y(ttmp116),.A(g166),.B(g2095));
AND2X1 AND_tmp117 (.Y(ttmp117),.A(g2078),.B(ttmp116));
AND2X1 AND_tmp118 (.Y(I5887),.A(g2083),.B(ttmp117));
AND2X1 AND2_1104 (.Y(g7823),.A(g1923),.B(g7479));
AND2X1 AND2_1105 (.Y(g4069),.A(g1762),.B(g2802));
AND2X1 AND_tmp119 (.Y(ttmp119),.A(g3015),.B(g11492));
AND2X1 AND_tmp120 (.Y(g11519),.A(g1317),.B(ttmp119));
AND2X1 AND2_1106 (.Y(g11176),.A(g506),.B(g11112));
AND2X1 AND2_1107 (.Y(g11092),.A(g837),.B(g10950));
AND2X1 AND2_1108 (.Y(g11154),.A(g330),.B(g10932));
AND2X1 AND2_1109 (.Y(g9608),.A(g7),.B(g9292));
AND2X1 AND2_1110 (.Y(g11637),.A(g11626),.B(g5446));
AND2X1 AND2_1111 (.Y(g2091),.A(g976),.B(g971));
AND2X1 AND2_1112 (.Y(g8406),.A(g695),.B(g8131));
AND2X1 AND2_1113 (.Y(g5254),.A(g4335),.B(g4165));
AND2X1 AND2_1114 (.Y(g7260),.A(g6752),.B(g2345));
AND2X1 AND2_1115 (.Y(g5150),.A(g1275),.B(g4678));
AND2X1 AND2_1116 (.Y(g8766),.A(g8612),.B(g5151));
AND2X1 AND2_1117 (.Y(g9588),.A(g3272),.B(g9173));
AND2X1 AND2_1118 (.Y(g8801),.A(g8742),.B(g8729));
AND2X1 AND2_1119 (.Y(g7063),.A(g5903),.B(g6582));
AND2X1 AND2_1120 (.Y(g10303),.A(g10208),.B(g9076));
AND2X1 AND2_1121 (.Y(g5009),.A(g1486),.B(g4640));
AND2X1 AND2_1122 (.Y(g9665),.A(g1314),.B(g9151));
AND2X1 AND2_1123 (.Y(g8748),.A(g7670),.B(g8656));
AND2X1 AND2_1124 (.Y(g11215),.A(g953),.B(g11160));
AND2X1 AND2_1125 (.Y(g10750),.A(g10687),.B(g3586));
AND2X1 AND_tmp121 (.Y(ttmp121),.A(g4921),.B(g3818));
AND2X1 AND_tmp122 (.Y(g5769),.A(g2112),.B(ttmp121));
AND2X1 AND2_1126 (.Y(g8755),.A(g7426),.B(g8671));
AND2X1 AND2_1127 (.Y(g6673),.A(g5305),.B(g5822));
AND2X1 AND2_1128 (.Y(g5212),.A(g1255),.B(g4726));
AND2X1 AND2_1129 (.Y(g7720),.A(g727),.B(g7232));
AND2X1 AND_tmp123 (.Y(ttmp123),.A(g5292),.B(g4609));
AND2X1 AND_tmp124 (.Y(g5918),.A(g2965),.B(ttmp123));
AND2X1 AND2_1130 (.Y(g8045),.A(g7547),.B(g5128));
AND2X1 AND2_1131 (.Y(g8173),.A(g7971),.B(g3112));
AND2X1 AND2_1132 (.Y(g11349),.A(g11288),.B(g7964));
AND2X1 AND2_1133 (.Y(g7843),.A(g7599),.B(g5919));
AND2X1 AND2_1134 (.Y(g9696),.A(g281),.B(g9432));
AND2X1 AND2_1135 (.Y(g6772),.A(g6228),.B(g722));
AND2X1 AND2_1136 (.Y(g6058),.A(g1035),.B(g5320));
AND2X1 AND2_1137 (.Y(g6531),.A(g79),.B(g6056));
AND2X1 AND2_1138 (.Y(g6743),.A(g4106),.B(g6146));
AND2X1 AND2_1139 (.Y(g6890),.A(g6752),.B(g6568));
AND2X1 AND2_1140 (.Y(g7549),.A(g7269),.B(g3829));
AND2X1 AND2_1141 (.Y(g8169),.A(g5265),.B(g7853));
AND2X1 AND2_1142 (.Y(g11304),.A(g5520),.B(g11245));
AND2X1 AND2_1143 (.Y(g9944),.A(g9924),.B(g9392));
AND2X1 AND2_1144 (.Y(g9240),.A(g6454),.B(g8962));
AND2X1 AND2_1145 (.Y(g8059),.A(g7592),.B(g5919));
AND2X1 AND2_1146 (.Y(g8718),.A(g8600),.B(g7903));
AND2X1 AND2_1147 (.Y(g8767),.A(g8616),.B(g5151));
AND2X1 AND2_1148 (.Y(g9316),.A(g8877),.B(g5708));
AND2X1 AND2_1149 (.Y(g7625),.A(g673),.B(g7085));
AND2X1 AND2_1150 (.Y(g8793),.A(g8644),.B(g8723));
AND2X1 AND2_1151 (.Y(g2940),.A(g2424),.B(g1654));
AND2X1 AND2_1152 (.Y(g4114),.A(g1351),.B(g3301));
AND2X1 AND2_1153 (.Y(g11636),.A(g11624),.B(g7936));
AND2X1 AND2_1154 (.Y(g10949),.A(g2947),.B(g10809));
AND2X1 AND2_1155 (.Y(g4870),.A(g237),.B(g3946));
AND2X1 AND2_1156 (.Y(g3563),.A(g3275),.B(g2126));
AND2X1 AND2_1157 (.Y(g10948),.A(g2223),.B(g10809));
AND2X1 AND2_1158 (.Y(g8246),.A(g7846),.B(g7442));
AND2X1 AND2_1159 (.Y(g5788),.A(g1540),.B(g5231));
AND2X1 AND2_1160 (.Y(g4008),.A(g2689),.B(g2276));
AND2X1 AND2_1161 (.Y(g9596),.A(g2649),.B(g9010));
AND2X1 AND2_1162 (.Y(g5249),.A(g1089),.B(g4747));
AND2X1 AND2_1163 (.Y(g11585),.A(g1321),.B(g11543));
AND2X1 AND2_1164 (.Y(g3089),.A(g2054),.B(g2050));
AND2X1 AND2_1165 (.Y(g4972),.A(g1436),.B(g4682));
AND2X1 AND2_1166 (.Y(g11554),.A(g2689),.B(g11519));
AND2X1 AND2_1167 (.Y(g7586),.A(g7096),.B(g5423));
AND2X1 AND2_1168 (.Y(g10673),.A(g10580),.B(g9450));
AND2X1 AND_tmp125 (.Y(ttmp125),.A(g3992),.B(g2493));
AND2X1 AND_tmp126 (.Y(g4806),.A(g3215),.B(ttmp125));
AND2X1 AND2_1169 (.Y(g5485),.A(g1914),.B(g4257));
AND2X1 AND2_1170 (.Y(g9936),.A(g9915),.B(g9624));
AND2X1 AND2_1171 (.Y(g2910),.A(g2424),.B(g1660));
AND2X1 AND2_1172 (.Y(g9317),.A(g6109),.B(g8875));
AND2X1 AND2_1173 (.Y(g10933),.A(g10853),.B(g3982));
AND2X1 AND2_1174 (.Y(g8388),.A(g8177),.B(g7689));
AND2X1 AND2_1175 (.Y(g4465),.A(g1117),.B(g3828));
AND2X1 AND2_1176 (.Y(g7141),.A(g6073),.B(g6716));
AND2X1 AND2_1177 (.Y(g10508),.A(g10391),.B(g2135));
AND2X1 AND2_1178 (.Y(g4230),.A(g1095),.B(g3638));
AND2X1 AND2_1179 (.Y(g10634),.A(g10604),.B(g3829));
AND2X1 AND2_1180 (.Y(g9601),.A(g922),.B(g9192));
AND2X1 AND2_1181 (.Y(g6126),.A(g5639),.B(g4319));
AND2X1 AND2_1182 (.Y(g6326),.A(g1250),.B(g5949));
AND2X1 AND2_1183 (.Y(g7710),.A(g700),.B(g7214));
AND2X1 AND2_1184 (.Y(g8028),.A(g7375),.B(g7436));
AND2X1 AND2_1185 (.Y(g6760),.A(g786),.B(g6221));
AND2X1 AND2_1186 (.Y(g5640),.A(g1059),.B(g4427));
AND2X1 AND2_1187 (.Y(g5031),.A(g1478),.B(g4640));
AND2X1 AND2_1188 (.Y(g4550),.A(g342),.B(g3586));
AND2X1 AND2_1189 (.Y(g7879),.A(g7610),.B(g3798));
AND2X1 AND2_1190 (.Y(g7962),.A(g7730),.B(g6712));
AND2X1 AND2_1191 (.Y(g9597),.A(g1170),.B(g9125));
AND2X1 AND2_1192 (.Y(g10452),.A(g10439),.B(g3388));
AND2X1 AND2_1193 (.Y(g4891),.A(g631),.B(g4739));
AND2X1 AND2_1194 (.Y(g5005),.A(g1490),.B(g4640));
AND2X1 AND2_1195 (.Y(g6423),.A(g4348),.B(g5784));
AND2X1 AND2_1196 (.Y(g8108),.A(g1891),.B(g7938));
AND2X1 AND_tmp127 (.Y(ttmp127),.A(g1289),.B(g3937));
AND2X1 AND_tmp128 (.Y(g4807),.A(g3015),.B(ttmp127));
AND2X1 AND2_1197 (.Y(g5911),.A(g3322),.B(g4977));
AND2X1 AND2_1198 (.Y(g9937),.A(g9916),.B(g9624));
AND2X1 AND2_1199 (.Y(g9840),.A(g9704),.B(g9747));
AND2X1 AND2_1200 (.Y(g10780),.A(g10723),.B(g5124));
AND2X1 AND2_1201 (.Y(g8217),.A(g1872),.B(g7883));
AND2X1 AND2_1202 (.Y(g11013),.A(g5209),.B(g10827));
AND2X1 AND2_1203 (.Y(g9390),.A(g1333),.B(g9151));
AND2X1 AND2_1204 (.Y(g11214),.A(g950),.B(g11159));
AND2X1 AND2_1205 (.Y(g6327),.A(g1255),.B(g5949));
AND2X1 AND2_1206 (.Y(g4342),.A(g1149),.B(g3719));
AND2X1 AND2_1207 (.Y(g5796),.A(g1564),.B(g5252));
AND2X1 AND2_1208 (.Y(g5473),.A(g4268),.B(g3518));
AND2X1 AND2_1209 (.Y(g6346),.A(g5038),.B(g5883));
AND2X1 AND2_1210 (.Y(g6633),.A(g354),.B(g6191));
AND2X1 AND2_1211 (.Y(g11005),.A(g5119),.B(g10827));
AND2X1 AND2_1212 (.Y(g8365),.A(g668),.B(g8240));
AND2X1 AND2_1213 (.Y(g8048),.A(g7558),.B(g5919));
AND2X1 AND2_1214 (.Y(g4481),.A(g1713),.B(g3906));
AND2X1 AND2_1215 (.Y(g4097),.A(g2677),.B(g2989));
AND2X1 AND2_1216 (.Y(g8055),.A(g7588),.B(g5128));
AND2X1 AND2_1217 (.Y(g4497),.A(g351),.B(g3586));
AND2X1 AND2_1218 (.Y(g9942),.A(g9922),.B(g9367));
AND2X1 AND2_1219 (.Y(g6696),.A(g5504),.B(g5850));
AND2X1 AND_tmp129 (.Y(ttmp129),.A(g1850),.B(g10665));
AND2X1 AND_tmp130 (.Y(g10731),.A(g5118),.B(ttmp129));
AND2X1 AND2_1220 (.Y(g8827),.A(g8552),.B(g8696));
AND2X1 AND2_1221 (.Y(g5540),.A(g1727),.B(g4315));
AND2X1 AND2_1222 (.Y(g4960),.A(g1403),.B(g4682));
AND2X1 AND2_1223 (.Y(g8846),.A(g8615),.B(g8712));
AND2X1 AND2_1224 (.Y(g6508),.A(g5983),.B(g3096));
AND2X1 AND2_1225 (.Y(g6240),.A(g182),.B(g5361));
AND2X1 AND2_1226 (.Y(g7931),.A(g2809),.B(g7446));
AND2X1 AND2_1227 (.Y(g5287),.A(g3876),.B(g4782));
AND2X1 AND2_1228 (.Y(g6472),.A(g5853),.B(g1936));
AND2X1 AND2_1229 (.Y(g11100),.A(g853),.B(g10950));
AND2X1 AND2_1230 (.Y(g11235),.A(g5443),.B(g11107));
AND2X1 AND2_1231 (.Y(g5199),.A(g1068),.B(g4719));
AND2X1 AND2_1232 (.Y(g6316),.A(g1270),.B(g5949));
AND2X1 AND2_1233 (.Y(g7515),.A(g7148),.B(g2855));
AND2X1 AND2_1234 (.Y(g10583),.A(g10518),.B(g10515));
AND2X1 AND2_1235 (.Y(g5781),.A(g1537),.B(g5222));
AND2X1 AND2_1236 (.Y(g8018),.A(g7742),.B(g7425));
AND2X1 AND2_1237 (.Y(g4401),.A(g2971),.B(g3772));
AND2X1 AND_tmp131 (.Y(ttmp131),.A(g6778),.B(g8925));
AND2X1 AND_tmp132 (.Y(g8994),.A(g8110),.B(ttmp131));
AND2X1 AND2_1238 (.Y(g2950),.A(g2424),.B(g1666));
AND2X1 AND2_1239 (.Y(g5510),.A(g1630),.B(g4280));
AND2X1 AND2_1240 (.Y(g6347),.A(g275),.B(g5890));
AND2X1 AND2_1241 (.Y(g9357),.A(g962),.B(g9223));
AND2X1 AND2_1242 (.Y(g4828),.A(g4106),.B(g695));
AND2X1 AND2_1243 (.Y(g11407),.A(g11339),.B(g5949));
AND2X1 AND2_1244 (.Y(g4727),.A(g386),.B(g3364));
AND2X1 AND2_1245 (.Y(g10357),.A(g10278),.B(g2462));
AND2X1 AND2_1246 (.Y(g10743),.A(g10639),.B(g4013));
AND2X1 AND2_1247 (.Y(g5259),.A(g627),.B(g4739));
AND2X1 AND2_1248 (.Y(g5694),.A(g162),.B(g5361));
AND2X1 AND2_1249 (.Y(g10769),.A(g10652),.B(g4840));
AND2X1 AND2_1250 (.Y(g11584),.A(g1318),.B(g11542));
AND2X1 AND2_1251 (.Y(g4932),.A(g1065),.B(g4442));
AND2X1 AND2_1252 (.Y(g10768),.A(g10649),.B(g4840));
AND2X1 AND2_1253 (.Y(g6820),.A(g1362),.B(g6596));
AND2X1 AND2_1254 (.Y(g4068),.A(g2719),.B(g2276));
AND2X1 AND2_1255 (.Y(g6317),.A(g1304),.B(g5949));
AND2X1 AND2_1256 (.Y(g5215),.A(g4276),.B(g3400));
AND2X1 AND2_1257 (.Y(g4576),.A(g530),.B(g4049));
AND2X1 AND2_1258 (.Y(g4866),.A(g231),.B(g3946));
AND2X1 AND2_1259 (.Y(g6775),.A(g822),.B(g6231));
AND2X1 AND2_1260 (.Y(g3829),.A(g2028),.B(g2728));
AND2X1 AND2_1261 (.Y(g10662),.A(g8892),.B(g10571));
AND2X1 AND2_1262 (.Y(g8101),.A(g6208),.B(g7877));
AND2X1 AND2_1263 (.Y(g5825),.A(g3204),.B(g5318));
AND2X1 AND_tmp133 (.Y(ttmp133),.A(g2421),.B(g2435));
AND2X1 AND_tmp134 (.Y(ttmp134),.A(g2396),.B(ttmp133));
AND2X1 AND_tmp135 (.Y(I6310),.A(g2407),.B(ttmp134));
AND2X1 AND2_1264 (.Y(g7884),.A(g7457),.B(g7022));
AND2X1 AND2_1265 (.Y(g5008),.A(g1292),.B(g4507));
AND2X1 AND2_1266 (.Y(g3974),.A(g231),.B(g3164));
AND2X1 AND2_1267 (.Y(g9949),.A(g9929),.B(g9392));
AND2X1 AND2_1268 (.Y(g2531),.A(g658),.B(g668));
AND2X1 AND2_1269 (.Y(g9292),.A(g8878),.B(g5708));
AND2X1 AND2_1270 (.Y(g10778),.A(g1027),.B(g10729));
AND2X1 AND2_1271 (.Y(g8041),.A(g7524),.B(g5128));
AND2X1 AND2_1272 (.Y(g6079),.A(g1053),.B(g5320));
AND2X1 AND2_1273 (.Y(g7235),.A(g6663),.B(g6447));
AND2X1 AND2_1274 (.Y(g9603),.A(g1173),.B(g9125));
AND2X1 AND2_1275 (.Y(g6840),.A(g248),.B(g6596));
AND2X1 AND2_1276 (.Y(g9850),.A(g9726),.B(g9560));
AND2X1 AND2_1277 (.Y(g7988),.A(g1878),.B(g7379));
AND2X1 AND2_1278 (.Y(g5228),.A(g1086),.B(g4734));
AND2X1 AND2_1279 (.Y(g7134),.A(g5587),.B(g6354));
AND2X1 AND2_1280 (.Y(g5934),.A(g5215),.B(g1965));
AND2X1 AND2_1281 (.Y(g5230),.A(g1265),.B(g4735));
AND2X1 AND2_1282 (.Y(g8168),.A(g5262),.B(g7853));
AND2X1 AND2_1283 (.Y(g9583),.A(g886),.B(g8995));
AND2X1 AND2_1284 (.Y(g10672),.A(g10579),.B(g9449));
AND2X1 AND2_1285 (.Y(g3287),.A(g802),.B(g2534));
AND2X1 AND2_1286 (.Y(g8772),.A(g8627),.B(g5151));
AND2X1 AND2_1287 (.Y(g4893),.A(g635),.B(g4739));
AND2X1 AND2_1288 (.Y(g10331),.A(g10256),.B(g3307));
AND2X1 AND2_1289 (.Y(g8505),.A(g8309),.B(g4789));
AND2X1 AND2_1290 (.Y(g10449),.A(g10420),.B(g3345));
AND2X1 AND2_1291 (.Y(g11273),.A(g5638),.B(g11195));
AND2X1 AND2_1292 (.Y(g8734),.A(g8626),.B(g7923));
AND2X1 AND2_1293 (.Y(g5913),.A(g1041),.B(g5320));
AND2X1 AND2_1294 (.Y(g10448),.A(g10421),.B(g3335));
AND2X1 AND2_1295 (.Y(g6163),.A(g4572),.B(g5354));
AND2X1 AND2_1296 (.Y(g6363),.A(g284),.B(g5901));
AND2X1 AND2_1297 (.Y(g7202),.A(g6349),.B(g4329));
AND2X1 AND2_1298 (.Y(g11463),.A(g11432),.B(g5446));
AND2X1 AND2_1299 (.Y(g8074),.A(g718),.B(g7826));
AND2X1 AND2_1300 (.Y(g4325),.A(g1166),.B(g3682));
AND2X1 AND2_1301 (.Y(g8474),.A(g8383),.B(g5285));
AND2X1 AND2_1302 (.Y(g11234),.A(g5424),.B(g11106));
AND2X1 AND2_1303 (.Y(g5266),.A(g718),.B(g4766));
AND2X1 AND2_1304 (.Y(g4483),.A(g336),.B(g3586));
AND2X1 AND2_1305 (.Y(g5248),.A(g673),.B(g4738));
AND2X1 AND2_1306 (.Y(g11514),.A(g11491),.B(g5151));
AND2X1 AND2_1307 (.Y(g5255),.A(g682),.B(g4754));
AND2X1 AND2_1308 (.Y(g4106),.A(g3284),.B(g686));
AND2X1 AND2_1309 (.Y(g2760),.A(g981),.B(g2091));
AND2X1 AND2_1310 (.Y(g5097),.A(g1786),.B(g4603));
AND2X1 AND2_1311 (.Y(g5726),.A(g1601),.B(g5167));
AND2X1 AND2_1312 (.Y(g5497),.A(g4296),.B(g3522));
AND2X1 AND2_1313 (.Y(g5354),.A(g2733),.B(g4460));
AND2X1 AND2_1314 (.Y(g7933),.A(g2814),.B(g7450));
AND2X1 AND2_1315 (.Y(g9617),.A(g9),.B(g9274));
AND2X1 AND2_1316 (.Y(g9906),.A(g9873),.B(g9683));
AND2X1 AND2_1317 (.Y(g11012),.A(g5196),.B(g10827));
AND2X1 AND2_1318 (.Y(g7050),.A(g5896),.B(g6575));
AND2X1 AND2_1319 (.Y(g10971),.A(g10849),.B(g3161));
AND2X1 AND2_1320 (.Y(g4904),.A(g1850),.B(g4243));
AND2X1 AND2_1321 (.Y(g10369),.A(g10361),.B(g3382));
AND2X1 AND2_1322 (.Y(g8400),.A(g6097),.B(g8234));
AND2X1 AND2_1323 (.Y(g4345),.A(g1169),.B(g3730));
AND2X1 AND2_1324 (.Y(g2161),.A(I5084),.B(I5085));
AND2X1 AND2_1325 (.Y(g5001),.A(g1300),.B(g4491));
AND2X1 AND2_1326 (.Y(g9945),.A(g9925),.B(g9392));
AND2X1 AND2_1327 (.Y(g7271),.A(g5028),.B(g6499));
AND2X1 AND2_1328 (.Y(g9709),.A(g1524),.B(g9490));
AND2X1 AND2_1329 (.Y(g4223),.A(g1003),.B(g3914));
AND2X1 AND2_1330 (.Y(g10716),.A(g10497),.B(g10675));
AND2X1 AND2_1331 (.Y(g11291),.A(g11247),.B(g4233));
AND2X1 AND2_1332 (.Y(g6661),.A(g73),.B(g6219));
AND2X1 AND2_1333 (.Y(g11173),.A(g491),.B(g11112));
AND2X1 AND2_1334 (.Y(g6075),.A(g549),.B(g5613));
AND2X1 AND2_1335 (.Y(g8023),.A(g7367),.B(g7430));
AND2X1 AND2_1336 (.Y(g9907),.A(g9888),.B(g9686));
AND2X1 AND2_1337 (.Y(g10582),.A(g10532),.B(g9473));
AND2X1 AND2_1338 (.Y(g5746),.A(g1589),.B(g5193));
AND2X1 AND2_1339 (.Y(g5221),.A(g1260),.B(g4730));
AND2X1 AND2_1340 (.Y(g9959),.A(g9950),.B(g9536));
AND2X1 AND2_1341 (.Y(g7674),.A(g7004),.B(g3880));
AND2X1 AND2_1342 (.Y(g9690),.A(g266),.B(g9432));
AND2X1 AND2_1343 (.Y(g6627),.A(g58),.B(g6181));
AND2X1 AND2_1344 (.Y(g5703),.A(g174),.B(g5361));
AND2X1 AND2_1345 (.Y(g4522),.A(g360),.B(g3586));
AND2X1 AND2_1346 (.Y(g4115),.A(g2689),.B(g3009));
AND2X1 AND2_1347 (.Y(g7541),.A(g7075),.B(g3109));
AND2X1 AND2_1348 (.Y(g10627),.A(g10548),.B(g4564));
AND2X1 AND2_1349 (.Y(g4047),.A(g2695),.B(g2276));
AND2X1 AND2_1350 (.Y(g6526),.A(g76),.B(g6052));
AND2X1 AND2_1351 (.Y(g2944),.A(g2424),.B(g1669));
AND2X1 AND2_1352 (.Y(g6646),.A(g360),.B(g6203));
AND2X1 AND2_1353 (.Y(g7132),.A(g6048),.B(g6702));
AND2X1 AND2_1354 (.Y(g11029),.A(g401),.B(g10974));
AND2X1 AND2_1355 (.Y(g8051),.A(g7572),.B(g5128));
AND2X1 AND2_1356 (.Y(g8127),.A(g1927),.B(g7949));
AND2X1 AND2_1357 (.Y(g7209),.A(g3804),.B(g6425));
AND2X1 AND2_1358 (.Y(g11028),.A(g396),.B(g10974));
AND2X1 AND2_1359 (.Y(g6439),.A(g4479),.B(g5919));
AND2X1 AND2_1360 (.Y(g10742),.A(g10655),.B(g3586));
AND2X1 AND2_1361 (.Y(g9110),.A(g8880),.B(g4790));
AND2X1 AND2_1362 (.Y(g10681),.A(g10567),.B(g3586));
AND2X1 AND2_1363 (.Y(g4537),.A(g444),.B(g3988));
AND2X1 AND2_1364 (.Y(g9663),.A(g959),.B(g9223));
AND2X1 AND2_1365 (.Y(g5349),.A(g2126),.B(g4617));
AND2X1 AND2_1366 (.Y(g8732),.A(g8624),.B(g7919));
AND2X1 AND2_1367 (.Y(g3807),.A(g3003),.B(g3062));
AND2X1 AND2_1368 (.Y(g8753),.A(g7414),.B(g8664));
AND2X1 AND2_1369 (.Y(g5848),.A(g3860),.B(g5519));
AND2X1 AND2_1370 (.Y(g8508),.A(g8411),.B(g7967));
AND2X1 AND2_1371 (.Y(g8072),.A(g700),.B(g7826));
AND2X1 AND2_1372 (.Y(g5699),.A(g1592),.B(g5117));
AND2X1 AND2_1373 (.Y(g11240),.A(g5481),.B(g11111));
AND2X1 AND2_1374 (.Y(g5398),.A(g4610),.B(g2224));
AND2X1 AND2_1375 (.Y(g6616),.A(g6105),.B(g3246));
AND2X1 AND2_1376 (.Y(g10690),.A(g10616),.B(g3863));
AND2X1 AND2_1377 (.Y(g8043),.A(g7582),.B(g5128));
AND2X1 AND2_1378 (.Y(g9590),.A(g895),.B(g8995));
AND2X1 AND2_1379 (.Y(g4128),.A(g1976),.B(g2779));
AND2X1 AND2_1380 (.Y(g6404),.A(g2132),.B(g5748));
AND2X1 AND2_1381 (.Y(g6647),.A(g5288),.B(g5808));
AND2X1 AND2_1382 (.Y(g10504),.A(g10389),.B(g2135));
AND2X1 AND2_1383 (.Y(g9657),.A(g919),.B(g9205));
AND2X1 AND2_1384 (.Y(g4542),.A(g366),.B(g3586));
AND2X1 AND2_1385 (.Y(g4330),.A(g1163),.B(g3693));
AND2X1 AND2_1386 (.Y(g3497),.A(g2804),.B(g1900));
AND2X1 AND2_1387 (.Y(g5524),.A(g1678),.B(g4291));
AND2X1 AND2_1388 (.Y(g8147),.A(g2955),.B(g7961));
AND2X1 AND2_1389 (.Y(g4554),.A(g542),.B(g3996));
AND2X1 AND2_1390 (.Y(g9899),.A(g9889),.B(g9367));
AND2X1 AND2_1391 (.Y(g5258),.A(g700),.B(g4756));
AND2X1 AND2_1392 (.Y(g7736),.A(g6951),.B(g3880));
AND2X1 AND2_1393 (.Y(g6224),.A(g1520),.B(g5151));
AND2X1 AND2_1394 (.Y(g10626),.A(g10547),.B(g4558));
AND2X1 AND2_1395 (.Y(g6320),.A(g1292),.B(g5949));
AND2X1 AND2_1396 (.Y(g7623),.A(g664),.B(g7079));
AND2X1 AND2_1397 (.Y(g10299),.A(g8892),.B(g10217));
AND2X1 AND2_1398 (.Y(g7889),.A(g7615),.B(g3814));
AND2X1 AND2_1399 (.Y(g10298),.A(g8892),.B(g10214));
AND2X1 AND2_1400 (.Y(g8413),.A(g722),.B(g8146));
AND2X1 AND2_1401 (.Y(g3979),.A(g237),.B(g3164));
AND2X1 AND2_1402 (.Y(g4902),.A(g1848),.B(g4243));
AND2X1 AND2_1403 (.Y(g5211),.A(g1080),.B(g4724));
AND2X1 AND2_1404 (.Y(g4512),.A(g357),.B(g3586));
AND2X1 AND2_1405 (.Y(g7722),.A(g7127),.B(g6449));
AND2X1 AND2_1406 (.Y(g9844),.A(g9714),.B(g9522));
AND2X1 AND2_1407 (.Y(g4490),.A(g1141),.B(g3913));
AND2X1 AND2_1408 (.Y(g4823),.A(g207),.B(g3946));
AND2X1 AND2_1409 (.Y(g6516),.A(g5993),.B(g3097));
AND2X1 AND2_1410 (.Y(g5026),.A(g1453),.B(g4640));
AND2X1 AND2_1411 (.Y(g8820),.A(g8705),.B(g5422));
AND2X1 AND2_1412 (.Y(g10737),.A(g10687),.B(g4840));
AND2X1 AND_tmp136 (.Y(ttmp136),.A(g6778),.B(g8849));
AND2X1 AND_tmp137 (.Y(g8936),.A(g8115),.B(ttmp136));
AND2X1 AND2_1413 (.Y(g10232),.A(g8892),.B(g10150));
AND2X1 AND2_1414 (.Y(g6771),.A(g263),.B(g5866));
AND2X1 AND2_1415 (.Y(g5170),.A(g1811),.B(g4680));
AND2X1 AND2_1416 (.Y(g8117),.A(g6236),.B(g7886));
AND2X1 AND2_1417 (.Y(g4529),.A(g448),.B(g3980));
AND2X1 AND2_1418 (.Y(g4348),.A(g3497),.B(g1909));
AND2X1 AND2_1419 (.Y(g9966),.A(g9956),.B(g9536));
AND2X1 AND2_1420 (.Y(g5280),.A(g4593),.B(g3052));
AND2X1 AND2_1421 (.Y(g7139),.A(g6060),.B(g6709));
AND2X1 AND2_1422 (.Y(g11099),.A(g382),.B(g10885));
AND2X1 AND2_1423 (.Y(g6892),.A(g6472),.B(g5805));
AND2X1 AND2_1424 (.Y(g9705),.A(g1580),.B(g9474));
AND2X1 AND2_1425 (.Y(g10512),.A(g10395),.B(g2135));
AND2X1 AND2_1426 (.Y(g11098),.A(g849),.B(g10950));
AND2X1 AND2_1427 (.Y(g8775),.A(g8628),.B(g5151));
AND2X1 AND2_1428 (.Y(g5083),.A(g3709),.B(g4586));
AND2X1 AND2_1429 (.Y(g5544),.A(g1687),.B(g4320));
AND2X1 AND2_1430 (.Y(g11272),.A(g5629),.B(g11193));
AND2X1 AND2_1431 (.Y(g5483),.A(g1621),.B(g4254));
AND2X1 AND2_1432 (.Y(g9948),.A(g9928),.B(g9392));
AND2X1 AND2_1433 (.Y(g4063),.A(g2713),.B(g2276));
AND2X1 AND2_1434 (.Y(g11462),.A(g11431),.B(g5446));
AND2X1 AND2_1435 (.Y(g6738),.A(g2531),.B(g6137));
AND2X1 AND2_1436 (.Y(g8060),.A(g7593),.B(g5919));
AND2X1 AND2_1437 (.Y(g6244),.A(g2255),.B(g5151));
AND2X1 AND2_1438 (.Y(g11032),.A(g416),.B(g10974));
AND2X1 AND2_1439 (.Y(g10445),.A(g10315),.B(g2135));
AND2X1 AND2_1440 (.Y(g9150),.A(g8882),.B(g4805));
AND2X1 AND2_1441 (.Y(g10316),.A(g10223),.B(g9097));
AND2X1 AND2_1442 (.Y(g5756),.A(g1531),.B(g5202));
AND2X1 AND2_1443 (.Y(g4720),.A(g1023),.B(g3914));
AND2X1 AND2_1444 (.Y(g9409),.A(g1721),.B(g9052));
AND2X1 AND2_1445 (.Y(g8995),.A(g6454),.B(g8929));
AND2X1 AND2_1446 (.Y(g6876),.A(g4070),.B(g6560));
AND2X1 AND2_1447 (.Y(g4989),.A(g1424),.B(g4682));
AND2X1 AND2_1448 (.Y(g9836),.A(g9737),.B(g9785));
AND2X1 AND_tmp138 (.Y(ttmp138),.A(g6061),.B(g4631));
AND2X1 AND_tmp139 (.Y(g6656),.A(g2733),.B(ttmp138));
AND2X1 AND2_1449 (.Y(g5514),.A(g1941),.B(g4284));
AND2X1 AND2_1450 (.Y(g8390),.A(g8268),.B(g6465));
AND2X1 AND2_1451 (.Y(g5003),.A(g1466),.B(g4640));
AND2X1 AND2_1452 (.Y(g9967),.A(g9957),.B(g9536));
AND2X1 AND2_1453 (.Y(g5145),.A(g1639),.B(g4673));
AND2X1 AND2_1454 (.Y(g4834),.A(g219),.B(g3946));
AND2X1 AND2_1455 (.Y(g4971),.A(g1419),.B(g4682));
AND2X1 AND2_1456 (.Y(g10753),.A(g10649),.B(g4013));
AND2X1 AND2_1457 (.Y(g5695),.A(g166),.B(g5361));
AND2X1 AND2_1458 (.Y(g7613),.A(g6940),.B(g5984));
AND2X1 AND2_1459 (.Y(g10736),.A(g10658),.B(g4840));
AND2X1 AND2_1460 (.Y(g11220),.A(g962),.B(g11054));
AND2X1 AND2_1461 (.Y(g7444),.A(g7277),.B(g5827));
AND2X1 AND2_1462 (.Y(g5536),.A(g4867),.B(g4298));
AND2X1 AND2_1463 (.Y(g6663),.A(g6064),.B(g2237));
AND2X1 AND2_1464 (.Y(g4670),.A(g192),.B(g3946));
AND2X1 AND2_1465 (.Y(g6824),.A(g1371),.B(g6596));
AND2X1 AND2_1466 (.Y(g4253),.A(g1074),.B(g3638));
AND2X1 AND2_1467 (.Y(g8250),.A(g2771),.B(g7907));
AND2X1 AND2_1468 (.Y(g8163),.A(g7960),.B(g3737));
AND2X1 AND2_1469 (.Y(g10764),.A(g10643),.B(g4840));
AND2X1 AND2_1470 (.Y(g5757),.A(g1552),.B(g5203));
AND2X1 AND2_1471 (.Y(g10365),.A(g10319),.B(g2135));
AND2X1 AND2_1472 (.Y(g8032),.A(g7385),.B(g7438));
AND2X1 AND2_1473 (.Y(g11591),.A(g2988),.B(g11561));
AND2X1 AND2_1474 (.Y(g8053),.A(g7583),.B(g5919));
AND2X1 AND2_1475 (.Y(g11147),.A(g321),.B(g10929));
AND2X1 AND2_1476 (.Y(g5522),.A(g1633),.B(g4289));
AND2X1 AND2_1477 (.Y(g5115),.A(g1394),.B(g4572));
AND2X1 AND2_1478 (.Y(g9837),.A(g9697),.B(g9751));
AND2X1 AND2_1479 (.Y(g9620),.A(g2653),.B(g9240));
AND2X1 AND2_1480 (.Y(g11151),.A(g327),.B(g10931));
AND2X1 AND2_1481 (.Y(g11172),.A(g486),.B(g11112));
AND2X1 AND2_1482 (.Y(g7885),.A(g7614),.B(g3812));
AND2X1 AND2_1483 (.Y(g6064),.A(g5398),.B(g2230));
AND2X1 AND_tmp140 (.Y(ttmp140),.A(g6368),.B(g8828));
AND2X1 AND_tmp141 (.Y(g8929),.A(g8095),.B(ttmp140));
AND2X1 AND2_1484 (.Y(g5595),.A(g1621),.B(g4524));
AND2X1 AND2_1485 (.Y(g5537),.A(g4143),.B(g4299));
AND2X1 AND2_1486 (.Y(g9842),.A(g9708),.B(g9516));
AND2X1 AND2_1487 (.Y(g4141),.A(g2707),.B(g3051));
AND2X1 AND2_1488 (.Y(g4341),.A(g339),.B(g3586));
AND2X1 AND2_1489 (.Y(g9192),.A(g6454),.B(g8955));
AND2X1 AND2_1490 (.Y(g7679),.A(g1950),.B(g6863));
AND2X1 AND2_1491 (.Y(g7378),.A(g6990),.B(g3880));
AND2X1 AND2_1492 (.Y(g5612),.A(g1627),.B(g4543));
AND2X1 AND2_1493 (.Y(g3939),.A(g213),.B(g3164));
AND2X1 AND2_1494 (.Y(g7135),.A(g869),.B(g6355));
AND2X1 AND2_1495 (.Y(g10970),.A(g10852),.B(g3390));
AND2X1 AND2_1496 (.Y(g11025),.A(g426),.B(g10974));
AND2X1 AND2_1497 (.Y(g9854),.A(g9730),.B(g9566));
AND2X1 AND2_1498 (.Y(g7182),.A(g1878),.B(g6720));
AND2X1 AND2_1499 (.Y(g9941),.A(g9921),.B(g9367));
AND2X1 AND2_1500 (.Y(g6194),.A(g554),.B(g5043));
AND2X1 AND2_1501 (.Y(g5128),.A(g4474),.B(g2733));
AND2X1 AND2_1502 (.Y(g4962),.A(g1651),.B(g4461));
AND2X1 AND2_1503 (.Y(g4358),.A(g1209),.B(g3747));
AND2X1 AND2_1504 (.Y(g8683),.A(g4803),.B(g8549));
AND2X1 AND2_1505 (.Y(g4506),.A(g1113),.B(g3944));
AND2X1 AND2_1506 (.Y(g6471),.A(g5224),.B(g6014));
AND2X1 AND2_1507 (.Y(g8778),.A(g8688),.B(g2317));
AND2X1 AND2_1508 (.Y(g11281),.A(g4948),.B(g11202));
AND2X1 AND2_1509 (.Y(g8735),.A(g7600),.B(g8632));
AND2X1 AND2_1510 (.Y(g11146),.A(g318),.B(g10928));
AND2X1 AND2_1511 (.Y(g3904),.A(g2948),.B(g2779));
AND2X1 AND2_1512 (.Y(g8075),.A(g727),.B(g7826));
AND2X1 AND2_1513 (.Y(g9829),.A(g9723),.B(g9785));
AND2X1 AND_tmp142 (.Y(ttmp142),.A(g6368),.B(g8828));
AND2X1 AND_tmp143 (.Y(g8949),.A(g8255),.B(ttmp142));
AND2X1 AND2_1514 (.Y(g7632),.A(g7184),.B(g5574));
AND2X1 AND2_1515 (.Y(g11290),.A(g11246),.B(g4226));
AND2X1 AND2_1516 (.Y(g6350),.A(g5837),.B(g4435));
AND2X1 AND2_1517 (.Y(g10599),.A(g10534),.B(g4365));
AND2X1 AND2_1518 (.Y(g5902),.A(g2555),.B(g4977));
AND2X1 AND_tmp144 (.Y(ttmp144),.A(g2407),.B(g2396));
AND2X1 AND_tmp145 (.Y(ttmp145),.A(g201),.B(ttmp144));
AND2X1 AND_tmp146 (.Y(I6337),.A(g2421),.B(ttmp145));
AND2X1 AND2_1519 (.Y(g2276),.A(g1765),.B(g1610));
AND2X1 AND2_1520 (.Y(g6438),.A(g5853),.B(g5797));
AND2X1 AND2_1521 (.Y(g5512),.A(g1660),.B(g4281));
AND2X1 AND2_1522 (.Y(g5090),.A(g1781),.B(g4592));
AND2X1 AND2_1523 (.Y(g7719),.A(g718),.B(g7227));
AND2X1 AND2_1524 (.Y(g2561),.A(g742),.B(g741));
AND2X1 AND2_1525 (.Y(g3695),.A(g1712),.B(g3015));
AND2X1 AND2_1526 (.Y(g8603),.A(g3983),.B(g8548));
AND2X1 AND2_1527 (.Y(g8039),.A(g7587),.B(g5128));
AND2X1 AND2_1528 (.Y(g9610),.A(g925),.B(g9192));
AND2X1 AND2_1529 (.Y(g3536),.A(g2390),.B(g3103));
AND2X1 AND2_1530 (.Y(g5529),.A(g4129),.B(g4288));
AND2X1 AND2_1531 (.Y(g5148),.A(g3088),.B(g4671));
AND2X1 AND2_1532 (.Y(g9124),.A(g8881),.B(g4802));
AND2X1 AND2_1533 (.Y(g9324),.A(g8879),.B(g5708));
AND2X1 AND2_1534 (.Y(g4559),.A(g2034),.B(g3829));
AND2X1 AND2_1535 (.Y(g10561),.A(g10549),.B(g4583));
AND2X1 AND2_1536 (.Y(g5698),.A(g1571),.B(g5116));
AND2X1 AND2_1537 (.Y(g11226),.A(g461),.B(g11057));
AND2X1 AND2_1538 (.Y(g10295),.A(g8892),.B(g10208));
AND2X1 AND2_1539 (.Y(g5260),.A(g1092),.B(g4758));
AND2X1 AND2_1540 (.Y(g10680),.A(g10564),.B(g3586));
AND2X1 AND2_1541 (.Y(g6822),.A(g231),.B(g6596));
AND2X1 AND2_1542 (.Y(g4905),.A(g1853),.B(g4243));
AND2X1 AND2_1543 (.Y(g11551),.A(g11538),.B(g4013));
AND2X1 AND2_1544 (.Y(g3047),.A(g1227),.B(g2306));
AND2X1 AND2_1545 (.Y(g9849),.A(g293),.B(g9768));
AND2X1 AND2_1546 (.Y(g5279),.A(g1766),.B(g4783));
AND2X1 AND2_1547 (.Y(g8404),.A(g686),.B(g8129));
AND2X1 AND2_1548 (.Y(g5720),.A(g170),.B(g5361));
AND2X1 AND2_1549 (.Y(g5318),.A(g4401),.B(g1857));
AND2X1 AND2_1550 (.Y(g8764),.A(g7443),.B(g8684));
AND2X1 AND2_1551 (.Y(g11376),.A(g11318),.B(g4277));
AND2X1 AND2_1552 (.Y(g11297),.A(g5490),.B(g11242));
AND2X1 AND2_1553 (.Y(g9898),.A(g9887),.B(g9367));
OR2X1 OR2_0 (.Y(g6895),.A(g6776),.B(g4875));
OR2X1 OR2_1 (.Y(g7189),.A(g6632),.B(g6053));
OR2X1 OR2_2 (.Y(g9510),.A(g9125),.B(g9111));
OR2X1 OR2_3 (.Y(g7297),.A(g7132),.B(g6323));
OR2X1 OR2_4 (.Y(g9088),.A(g8927),.B(g8381));
OR2X1 OR2_5 (.Y(g9923),.A(g9865),.B(g9707));
OR2X1 OR2_6 (.Y(g6485),.A(g5848),.B(g5067));
OR2X1 OR2_7 (.Y(g8771),.A(g5483),.B(g8652));
OR2X1 OR2_8 (.Y(g5813),.A(g5617),.B(g4869));
OR2X1 OR2_9 (.Y(g7963),.A(g7687),.B(g7182));
OR2X1 OR2_10 (.Y(g10643),.A(g10624),.B(g7736));
OR2X1 OR_tmp147 (.Y(ttmp147),.A(g9592),.B(g9759));
OR2X1 OR_tmp148 (.Y(g9886),.A(g9607),.B(ttmp147));
OR2X1 OR_tmp149 (.Y(ttmp149),.A(g9899),.B(g9803));
OR2X1 OR_tmp150 (.Y(g9951),.A(g9902),.B(ttmp149));
OR2X1 OR2_11 (.Y(g11625),.A(g6535),.B(g11597));
OR2X1 OR2_12 (.Y(g8945),.A(g8801),.B(g8710));
OR2X1 OR2_13 (.Y(g10489),.A(g4961),.B(g10367));
OR2X1 OR2_14 (.Y(g10559),.A(g4141),.B(g10512));
OR2X1 OR2_15 (.Y(g10558),.A(g4126),.B(g10510));
OR2X1 OR2_16 (.Y(g11338),.A(g11283),.B(g11178));
OR2X1 OR2_17 (.Y(g8435),.A(g8403),.B(g8075));
OR2X1 OR2_18 (.Y(g10544),.A(g5511),.B(g10495));
OR2X1 OR2_19 (.Y(g6911),.A(g6342),.B(g5681));
OR2X1 OR2_20 (.Y(g10865),.A(g5538),.B(g10752));
OR2X1 OR2_21 (.Y(g3698),.A(g3121),.B(g2480));
OR2X1 OR2_22 (.Y(g8214),.A(g7472),.B(g8004));
OR2X1 OR2_23 (.Y(g6124),.A(g5181),.B(g5188));
OR2X1 OR2_24 (.Y(g6469),.A(g5698),.B(g4959));
OR2X1 OR2_25 (.Y(g5587),.A(g4714),.B(g3904));
OR2X1 OR2_26 (.Y(g6177),.A(g5444),.B(g4712));
OR2X1 OR_tmp151 (.Y(ttmp151),.A(g9205),.B(g9192));
OR2X1 OR_tmp152 (.Y(I14585),.A(g8995),.B(ttmp151));
OR2X1 OR2_27 (.Y(g9891),.A(g9741),.B(g9760));
OR2X1 OR2_28 (.Y(g9913),.A(g9849),.B(g9691));
OR2X1 OR_tmp153 (.Y(ttmp153),.A(g486),.B(g481));
OR2X1 OR_tmp154 (.Y(ttmp154),.A(g496),.B(ttmp153));
OR2X1 OR_tmp155 (.Y(I5600),.A(g491),.B(ttmp154));
OR2X1 OR2_29 (.Y(g11257),.A(g11234),.B(g11019));
OR2X1 OR2_30 (.Y(g8236),.A(g7526),.B(g8001));
OR2X1 OR2_31 (.Y(g7385),.A(g7235),.B(g6746));
OR2X1 OR2_32 (.Y(g6898),.A(g6790),.B(g4881));
OR2X1 OR2_33 (.Y(g6900),.A(g6787),.B(g6246));
OR2X1 OR2_34 (.Y(g4264),.A(g4048),.B(g4053));
OR2X1 OR_tmp156 (.Y(ttmp156),.A(g9420),.B(g9489));
OR2X1 OR_tmp157 (.Y(g9726),.A(g9411),.B(ttmp156));
OR2X1 OR2_35 (.Y(g6088),.A(g5260),.B(g4522));
OR2X1 OR2_36 (.Y(g6923),.A(g6353),.B(g5695));
OR2X1 OR2_37 (.Y(g8194),.A(g5168),.B(g7940));
OR2X1 OR_tmp158 (.Y(ttmp158),.A(g9292),.B(g9274));
OR2X1 OR_tmp159 (.Y(g9676),.A(g9454),.B(ttmp158));
OR2X1 OR2_38 (.Y(g11256),.A(g11186),.B(g11018));
OR2X1 OR2_39 (.Y(g3860),.A(g3107),.B(g2167));
OR2X1 OR2_40 (.Y(g11280),.A(g11254),.B(g11153));
OR2X1 OR_tmp160 (.Y(ttmp160),.A(g9362),.B(I14866));
OR2X1 OR_tmp161 (.Y(ttmp161),.A(g9650),.B(ttmp160));
OR2X1 OR_tmp162 (.Y(g9727),.A(g9663),.B(ttmp161));
OR2X1 OR2_41 (.Y(g4997),.A(g4581),.B(g4584));
OR2X1 OR2_42 (.Y(g11624),.A(g11595),.B(g11571));
OR2X1 OR2_43 (.Y(g11300),.A(g11213),.B(g11091));
OR2X1 OR2_44 (.Y(g4238),.A(g3999),.B(g4007));
OR2X1 OR2_45 (.Y(g8814),.A(g7945),.B(g8728));
OR2X1 OR2_46 (.Y(g10401),.A(g9317),.B(g10291));
OR2X1 OR2_47 (.Y(g8773),.A(g5491),.B(g8653));
OR2X1 OR2_48 (.Y(g11231),.A(g11156),.B(g11013));
OR2X1 OR2_49 (.Y(g10864),.A(g5532),.B(g10751));
OR2X1 OR2_50 (.Y(g9624),.A(g9316),.B(g9313));
OR2X1 OR_tmp163 (.Y(ttmp163),.A(g9939),.B(g9669));
OR2X1 OR_tmp164 (.Y(g9953),.A(g9945),.B(ttmp163));
OR2X1 OR2_51 (.Y(g6122),.A(g5172),.B(g5180));
OR2X1 OR2_52 (.Y(g6465),.A(g5825),.B(g5041));
OR2X1 OR2_53 (.Y(g6934),.A(g6363),.B(g5720));
OR2X1 OR2_54 (.Y(g7664),.A(g6855),.B(g4084));
OR2X1 OR2_55 (.Y(g7246),.A(g6465),.B(g6003));
OR2X1 OR2_56 (.Y(g7203),.A(g6640),.B(g6058));
OR2X1 OR2_57 (.Y(g6096),.A(g5268),.B(g4542));
OR2X1 OR2_58 (.Y(g9747),.A(g9173),.B(g9509));
OR2X1 OR2_59 (.Y(g11314),.A(g11224),.B(g11102));
OR2X1 OR2_60 (.Y(g10733),.A(g5227),.B(g10674));
OR2X1 OR2_61 (.Y(g8921),.A(g8827),.B(g8748));
OR2X1 OR_tmp165 (.Y(ttmp165),.A(g9624),.B(g9785));
OR2X1 OR_tmp166 (.Y(ttmp166),.A(g7853),.B(ttmp165));
OR2X1 OR_tmp167 (.Y(I15054),.A(g9782),.B(ttmp166));
OR2X1 OR2_62 (.Y(g11269),.A(g11196),.B(g11031));
OR2X1 OR2_63 (.Y(g5555),.A(g4389),.B(g4397));
OR2X1 OR2_64 (.Y(g11268),.A(g11194),.B(g11030));
OR2X1 OR2_65 (.Y(g10485),.A(g9317),.B(g10376));
OR2X1 OR2_66 (.Y(g10555),.A(g4103),.B(g10504));
OR2X1 OR2_67 (.Y(g6481),.A(g5722),.B(g4972));
OR2X1 OR2_68 (.Y(g10712),.A(g10662),.B(g9531));
OR2X1 OR2_69 (.Y(g11335),.A(g11279),.B(g11175));
OR2X1 OR2_70 (.Y(g8249),.A(g8018),.B(g7710));
OR2X1 OR2_71 (.Y(g7638),.A(g7265),.B(g6488));
OR2X1 OR2_72 (.Y(g10567),.A(g10514),.B(g7378));
OR2X1 OR2_73 (.Y(g11487),.A(g6662),.B(g11464));
OR2X1 OR_tmp168 (.Y(ttmp168),.A(g9852),.B(g9882));
OR2X1 OR_tmp169 (.Y(ttmp169),.A(g9839),.B(ttmp168));
OR2X1 OR_tmp170 (.Y(I15210),.A(g9964),.B(ttmp169));
OR2X1 OR_tmp171 (.Y(ttmp171),.A(g2096),.B(g2088));
OR2X1 OR_tmp172 (.Y(ttmp172),.A(g2102),.B(ttmp171));
OR2X1 OR_tmp173 (.Y(I5805),.A(g2099),.B(ttmp172));
OR2X1 OR2_74 (.Y(g8941),.A(g8796),.B(g8706));
OR2X1 OR2_75 (.Y(g11443),.A(g7130),.B(g11407));
OR2X1 OR2_76 (.Y(g4231),.A(g3991),.B(g3998));
OR2X1 OR2_77 (.Y(g11278),.A(g11253),.B(g11150));
OR2X1 OR_tmp174 (.Y(ttmp174),.A(g9624),.B(g9785));
OR2X1 OR_tmp175 (.Y(ttmp175),.A(g7853),.B(ttmp174));
OR2X1 OR_tmp176 (.Y(I15039),.A(g9809),.B(ttmp175));
OR2X1 OR2_78 (.Y(g11286),.A(g10670),.B(g11209));
OR2X1 OR2_79 (.Y(g8431),.A(g8387),.B(g8071));
OR2X1 OR2_80 (.Y(g7133),.A(g6616),.B(g3067));
OR2X1 OR2_81 (.Y(g11306),.A(g11216),.B(g11095));
OR2X1 OR2_82 (.Y(g8252),.A(g7988),.B(g7679));
OR2X1 OR2_83 (.Y(g8812),.A(g7939),.B(g8724));
OR2X1 OR2_84 (.Y(g7846),.A(g7722),.B(g7241));
OR2X1 OR2_85 (.Y(g3875),.A(g3275),.B(g12));
OR2X1 OR2_86 (.Y(g5996),.A(g5473),.B(g3908));
OR2X1 OR2_87 (.Y(g6592),.A(g5100),.B(g5882));
OR2X1 OR2_88 (.Y(g8286),.A(g8107),.B(g7823));
OR2X1 OR2_89 (.Y(g10501),.A(g4161),.B(g10445));
OR2X1 OR2_90 (.Y(g10728),.A(g4973),.B(g10642));
OR2X1 OR2_91 (.Y(g8270),.A(g7894),.B(g3434));
OR2X1 OR2_92 (.Y(g7290),.A(g7046),.B(g6316));
OR2X1 OR2_93 (.Y(g6068),.A(g5220),.B(g4497));
OR2X1 OR2_94 (.Y(g6468),.A(g5690),.B(g4950));
OR2X1 OR2_95 (.Y(g11217),.A(g11144),.B(g11005));
OR2X1 OR2_96 (.Y(g11478),.A(g6532),.B(g11455));
OR2X1 OR_tmp177 (.Y(ttmp177),.A(g9328),.B(g9324));
OR2X1 OR_tmp178 (.Y(ttmp178),.A(g9335),.B(ttmp177));
OR2X1 OR_tmp179 (.Y(g9536),.A(g9331),.B(ttmp178));
OR2X1 OR2_97 (.Y(g5981),.A(g5074),.B(g4383));
OR2X1 OR2_98 (.Y(g11486),.A(g6654),.B(g11463));
OR2X1 OR2_99 (.Y(g8377),.A(g8185),.B(g7958));
OR2X1 OR2_100 (.Y(g8206),.A(g7459),.B(g8007));
OR2X1 OR2_101 (.Y(g11580),.A(g11413),.B(g11544));
OR2X1 OR2_102 (.Y(g8287),.A(g8117),.B(g7824));
OR2X1 OR2_103 (.Y(g11223),.A(g11147),.B(g11008));
OR2X1 OR2_104 (.Y(g9522),.A(g9173),.B(g9125));
OR2X1 OR2_105 (.Y(g8199),.A(g7902),.B(g7444));
OR2X1 OR2_106 (.Y(g5802),.A(g5601),.B(g4837));
OR2X1 OR2_107 (.Y(g11321),.A(g11230),.B(g11105));
OR2X1 OR2_108 (.Y(g6524),.A(g5746),.B(g4996));
OR2X1 OR2_109 (.Y(g10664),.A(g10240),.B(g10582));
OR2X1 OR2_110 (.Y(g7257),.A(g6701),.B(g4725));
OR2X1 OR2_111 (.Y(g7301),.A(g7140),.B(g6327));
OR2X1 OR2_112 (.Y(g10484),.A(g9317),.B(g10400));
OR2X1 OR2_113 (.Y(g10554),.A(g4097),.B(g10503));
OR2X1 OR2_114 (.Y(g8259),.A(g8028),.B(g7719));
OR2X1 OR2_115 (.Y(g11334),.A(g11277),.B(g11174));
OR2X1 OR2_116 (.Y(g8819),.A(g7957),.B(g8734));
OR2X1 OR2_117 (.Y(g8923),.A(g8846),.B(g8763));
OR2X1 OR2_118 (.Y(g8488),.A(g3664),.B(g8390));
OR2X1 OR2_119 (.Y(g7441),.A(g7271),.B(g6789));
OR2X1 OR2_120 (.Y(g6026),.A(g5507),.B(g3970));
OR2X1 OR2_121 (.Y(g10799),.A(g6225),.B(g10769));
OR2X1 OR2_122 (.Y(g10798),.A(g6217),.B(g10768));
OR2X1 OR2_123 (.Y(g10805),.A(g10759),.B(g10760));
OR2X1 OR2_124 (.Y(g10732),.A(g4358),.B(g10661));
OR2X1 OR2_125 (.Y(g6061),.A(g5204),.B(g4));
OR2X1 OR2_126 (.Y(g9512),.A(g9151),.B(g9125));
OR2X1 OR2_127 (.Y(g10013),.A(I15214),.B(I15215));
OR2X1 OR2_128 (.Y(g8806),.A(g7931),.B(g8718));
OR2X1 OR2_129 (.Y(g8943),.A(g8837),.B(g8749));
OR2X1 OR2_130 (.Y(g11293),.A(g11211),.B(g10818));
OR2X1 OR2_131 (.Y(g11265),.A(g11189),.B(g11027));
OR2X1 OR2_132 (.Y(g8887),.A(g8842),.B(g8755));
OR2X1 OR2_133 (.Y(g5838),.A(g5612),.B(g4866));
OR2X1 OR2_134 (.Y(g6514),.A(g5738),.B(g4992));
OR2X1 OR2_135 (.Y(g8322),.A(g8136),.B(g6891));
OR2X1 OR2_136 (.Y(g8230),.A(g7515),.B(g7991));
OR2X1 OR2_137 (.Y(g5809),.A(g5611),.B(g4865));
OR2X1 OR2_138 (.Y(g8433),.A(g8399),.B(g8073));
OR2X1 OR2_139 (.Y(g11579),.A(g5123),.B(g11551));
OR2X1 OR2_140 (.Y(g10771),.A(g5533),.B(g10684));
OR2X1 OR2_141 (.Y(g11615),.A(g11601),.B(g11592));
OR2X1 OR2_142 (.Y(g9367),.A(g9335),.B(g9331));
OR2X1 OR_tmp180 (.Y(ttmp180),.A(g9594),.B(g9750));
OR2X1 OR_tmp181 (.Y(g9872),.A(g9617),.B(ttmp180));
OR2X1 OR2_143 (.Y(g6522),.A(g5744),.B(g4994));
OR2X1 OR2_144 (.Y(g8266),.A(g7885),.B(g3412));
OR2X1 OR2_145 (.Y(g10414),.A(g10300),.B(g9534));
OR2X1 OR2_146 (.Y(g11275),.A(g11248),.B(g11148));
OR2X1 OR2_147 (.Y(g11430),.A(g11387),.B(g4006));
OR2X1 OR2_148 (.Y(g8248),.A(g8014),.B(g7707));
OR2X1 OR_tmp182 (.Y(ttmp182),.A(g9292),.B(g9274));
OR2X1 OR_tmp183 (.Y(g9686),.A(g9454),.B(ttmp182));
OR2X1 OR2_149 (.Y(g8815),.A(g7948),.B(g8730));
OR2X1 OR2_150 (.Y(g7183),.A(g6623),.B(g6046));
OR2X1 OR2_151 (.Y(g5983),.A(g5084),.B(g4392));
OR2X1 OR2_152 (.Y(g8154),.A(g7891),.B(g6879));
OR2X1 OR2_153 (.Y(g6537),.A(g5781),.B(g5005));
OR2X1 OR2_154 (.Y(g4309),.A(g4069),.B(g4079));
OR2X1 OR2_155 (.Y(g10725),.A(g4962),.B(g10634));
OR2X1 OR2_156 (.Y(g6243),.A(g5537),.B(g4774));
OR2X1 OR_tmp184 (.Y(ttmp184),.A(g2380),.B(g2372));
OR2X1 OR_tmp185 (.Y(ttmp185),.A(g2405),.B(ttmp184));
OR2X1 OR_tmp186 (.Y(I6351),.A(g2389),.B(ttmp185));
OR2X1 OR_tmp187 (.Y(ttmp187),.A(g9151),.B(g9125));
OR2X1 OR_tmp188 (.Y(g9519),.A(g9173),.B(ttmp187));
OR2X1 OR2_157 (.Y(g9740),.A(g9418),.B(g9505));
OR2X1 OR2_158 (.Y(g8267),.A(g7889),.B(g3422));
OR2X1 OR_tmp189 (.Y(ttmp189),.A(g10668),.B(I16427));
OR2X1 OR_tmp190 (.Y(g10744),.A(g10600),.B(ttmp189));
OR2X1 OR2_159 (.Y(g6542),.A(g5789),.B(g5010));
OR2X1 OR2_160 (.Y(g7303),.A(g7145),.B(g6329));
OR2X1 OR2_161 (.Y(g10652),.A(g10627),.B(g7743));
OR2X1 OR2_162 (.Y(g5036),.A(g4871),.B(g4162));
OR2X1 OR2_163 (.Y(g7240),.A(g6687),.B(g6095));
OR2X1 OR2_164 (.Y(g8221),.A(g7496),.B(g7993));
OR2X1 OR2_165 (.Y(g6902),.A(g6794),.B(g4223));
OR2X1 OR_tmp191 (.Y(ttmp191),.A(g9205),.B(g9192));
OR2X1 OR_tmp192 (.Y(I14776),.A(g8995),.B(ttmp191));
OR2X1 OR2_166 (.Y(g10500),.A(g4157),.B(g10442));
OR2X1 OR2_167 (.Y(g4052),.A(g2862),.B(g2515));
OR2X1 OR_tmp193 (.Y(ttmp193),.A(g9610),.B(g9602));
OR2X1 OR_tmp194 (.Y(ttmp194),.A(g9585),.B(ttmp193));
OR2X1 OR_tmp195 (.Y(I14858),.A(g9595),.B(ttmp194));
OR2X1 OR2_168 (.Y(g6529),.A(g5757),.B(g5000));
OR2X1 OR2_169 (.Y(g11264),.A(g11188),.B(g11026));
OR2X1 OR_tmp196 (.Y(ttmp196),.A(g9934),.B(g9830));
OR2X1 OR_tmp197 (.Y(ttmp197),.A(g8169),.B(ttmp196));
OR2X1 OR_tmp198 (.Y(I15209),.A(g9905),.B(ttmp197));
OR2X1 OR2_170 (.Y(g8241),.A(g7536),.B(g7989));
OR2X1 OR2_171 (.Y(g10795),.A(g6199),.B(g10764));
OR2X1 OR2_172 (.Y(g11607),.A(g11586),.B(g11557));
OR2X1 OR2_173 (.Y(g8644),.A(g8123),.B(g8464));
OR2X1 OR_tmp199 (.Y(ttmp199),.A(g3348),.B(g1570));
OR2X1 OR_tmp200 (.Y(g4682),.A(g3563),.B(ttmp199));
OR2X1 OR2_174 (.Y(g8818),.A(g7955),.B(g8733));
OR2X1 OR2_175 (.Y(g2984),.A(g2528),.B(g2522));
OR2X1 OR2_176 (.Y(g9931),.A(g8931),.B(g9900));
OR2X1 OR2_177 (.Y(g3414),.A(g2911),.B(g2917));
OR2X1 OR2_178 (.Y(g9515),.A(g9173),.B(g9151));
OR2X1 OR2_179 (.Y(g10724),.A(g10312),.B(g10672));
OR2X1 OR2_180 (.Y(g7294),.A(g7068),.B(g6320));
OR2X1 OR2_181 (.Y(g5189),.A(g4345),.B(g3496));
OR2X1 OR2_182 (.Y(g8614),.A(g8365),.B(g8510));
OR2X1 OR2_183 (.Y(g3513),.A(g3118),.B(g2180));
OR2X1 OR2_184 (.Y(g6909),.A(g6346),.B(g5684));
OR2X1 OR_tmp201 (.Y(ttmp201),.A(g386),.B(g426));
OR2X1 OR_tmp202 (.Y(ttmp202),.A(g396),.B(ttmp201));
OR2X1 OR_tmp203 (.Y(I5571),.A(g391),.B(ttmp202));
OR2X1 OR2_185 (.Y(g4283),.A(g4059),.B(g4063));
OR2X1 OR2_186 (.Y(g8939),.A(g8791),.B(g8701));
OR2X1 OR2_187 (.Y(g2514),.A(I5599),.B(I5600));
OR2X1 OR2_188 (.Y(g11327),.A(g11297),.B(g11167));
OR2X1 OR2_189 (.Y(g8187),.A(g7542),.B(g7998));
OR2X1 OR2_190 (.Y(g11606),.A(g11585),.B(g11556));
OR2X1 OR2_191 (.Y(g11303),.A(g11214),.B(g11092));
OR2X1 OR2_192 (.Y(g5309),.A(g3664),.B(g4401));
OR2X1 OR_tmp204 (.Y(ttmp204),.A(g9125),.B(g9111));
OR2X1 OR_tmp205 (.Y(g9528),.A(g9151),.B(ttmp204));
OR2X1 OR2_193 (.Y(g8200),.A(g7535),.B(g8008));
OR2X1 OR_tmp206 (.Y(ttmp206),.A(g829),.B(I5629));
OR2X1 OR_tmp207 (.Y(g2522),.A(g833),.B(ttmp206));
OR2X1 OR_tmp208 (.Y(ttmp208),.A(g1113),.B(I5363));
OR2X1 OR_tmp209 (.Y(ttmp209),.A(g1163),.B(ttmp208));
OR2X1 OR_tmp210 (.Y(g2315),.A(g1166),.B(ttmp209));
OR2X1 OR2_194 (.Y(g6506),.A(g5731),.B(g4989));
OR2X1 OR2_195 (.Y(g10649),.A(g10626),.B(g7741));
OR2X1 OR2_196 (.Y(g8159),.A(g7895),.B(g6886));
OR2X1 OR2_197 (.Y(g7626),.A(g7060),.B(g5267));
OR2X1 OR2_198 (.Y(g10770),.A(g5525),.B(g10682));
OR2X1 OR2_199 (.Y(g9566),.A(g9052),.B(g9030));
OR2X1 OR2_200 (.Y(g11483),.A(g6633),.B(g11460));
OR2X1 OR2_201 (.Y(g8811),.A(g7935),.B(g8722));
OR2X1 OR_tmp211 (.Y(ttmp211),.A(g5205),.B(g8465));
OR2X1 OR_tmp212 (.Y(g8642),.A(g5236),.B(ttmp211));
OR2X1 OR2_202 (.Y(g6545),.A(g5795),.B(g5025));
OR2X1 OR2_203 (.Y(g10767),.A(g5500),.B(g10681));
OR2X1 OR2_204 (.Y(g11326),.A(g11296),.B(g11166));
OR2X1 OR2_205 (.Y(g10898),.A(g4220),.B(g10777));
OR2X1 OR2_206 (.Y(g11252),.A(g11099),.B(g10969));
OR2X1 OR2_207 (.Y(g10719),.A(g10303),.B(g10666));
OR2X1 OR2_208 (.Y(g4609),.A(g3400),.B(g119));
OR2X1 OR2_209 (.Y(g6507),.A(g5732),.B(g4990));
OR2X1 OR2_210 (.Y(g10718),.A(g6238),.B(g10706));
OR2X1 OR2_211 (.Y(g10521),.A(I16148),.B(I16149));
OR2X1 OR2_212 (.Y(g7075),.A(g5104),.B(g6530));
OR2X1 OR2_213 (.Y(g7292),.A(g7055),.B(g6318));
OR2X1 OR2_214 (.Y(g10861),.A(g5523),.B(g10745));
OR2X1 OR2_215 (.Y(g8417),.A(g8246),.B(g7721));
OR2X1 OR2_216 (.Y(g6515),.A(g5739),.B(g4993));
OR2X1 OR_tmp213 (.Y(ttmp213),.A(g9601),.B(g9596));
OR2X1 OR_tmp214 (.Y(ttmp214),.A(g9583),.B(ttmp213));
OR2X1 OR_tmp215 (.Y(I14855),.A(g9593),.B(ttmp214));
OR2X1 OR_tmp216 (.Y(ttmp216),.A(g9850),.B(g9878));
OR2X1 OR_tmp217 (.Y(ttmp217),.A(g9838),.B(ttmp216));
OR2X1 OR_tmp218 (.Y(I15205),.A(g9963),.B(ttmp217));
OR2X1 OR_tmp219 (.Y(ttmp219),.A(g9624),.B(g9785));
OR2X1 OR_tmp220 (.Y(ttmp220),.A(g7853),.B(ttmp219));
OR2X1 OR_tmp221 (.Y(I15051),.A(g9673),.B(ttmp220));
OR2X1 OR_tmp222 (.Y(ttmp222),.A(g9419),.B(g9615));
OR2X1 OR_tmp223 (.Y(g9724),.A(g9409),.B(ttmp222));
OR2X1 OR2_217 (.Y(g6528),.A(g5756),.B(g4999));
OR2X1 OR2_218 (.Y(g8823),.A(g8778),.B(g8693));
OR2X1 OR2_219 (.Y(g7503),.A(g6887),.B(g6430));
OR2X1 OR2_220 (.Y(g8148),.A(g7884),.B(g6872));
OR2X1 OR2_221 (.Y(g8649),.A(g8499),.B(g4519));
OR2X1 OR2_222 (.Y(g3584),.A(g2863),.B(g2516));
OR2X1 OR2_223 (.Y(g10776),.A(g5544),.B(g10758));
OR2X1 OR_tmp224 (.Y(ttmp224),.A(g9292),.B(g9274));
OR2X1 OR_tmp225 (.Y(g9680),.A(g9454),.B(ttmp224));
OR2X1 OR2_224 (.Y(g10859),.A(g5512),.B(g10742));
OR2X1 OR_tmp226 (.Y(ttmp226),.A(g9609),.B(g9619));
OR2X1 OR_tmp227 (.Y(I14866),.A(g9590),.B(ttmp226));
OR2X1 OR2_225 (.Y(g7299),.A(g7138),.B(g6325));
OR2X1 OR2_226 (.Y(g10858),.A(g5501),.B(g10741));
OR2X1 OR2_227 (.Y(g8193),.A(g5145),.B(g7937));
OR2X1 OR_tmp228 (.Y(ttmp228),.A(g9125),.B(g9111));
OR2X1 OR_tmp229 (.Y(g9511),.A(g9151),.B(ttmp228));
OR2X1 OR2_228 (.Y(g7738),.A(g7200),.B(g6738));
OR2X1 OR2_229 (.Y(g7244),.A(g6699),.B(g4720));
OR2X1 OR2_230 (.Y(g3425),.A(g2895),.B(g2910));
OR2X1 OR2_231 (.Y(g7478),.A(g6884),.B(g6423));
OR2X1 OR_tmp230 (.Y(ttmp230),.A(g9366),.B(g9654));
OR2X1 OR_tmp231 (.Y(g9714),.A(g9664),.B(ttmp230));
OR2X1 OR2_232 (.Y(g10025),.A(I15224),.B(I15225));
OR2X1 OR2_233 (.Y(g6908),.A(g6345),.B(g4229));
OR2X1 OR2_234 (.Y(g5028),.A(g4836),.B(g4128));
OR2X1 OR2_235 (.Y(g8253),.A(g8023),.B(g7718));
OR2X1 OR2_236 (.Y(g8938),.A(g8789),.B(g8699));
OR2X1 OR2_237 (.Y(g8813),.A(g7943),.B(g8726));
OR2X1 OR2_238 (.Y(g9736),.A(g9430),.B(g9416));
OR2X1 OR2_239 (.Y(g9968),.A(I15171),.B(I15172));
OR2X1 OR2_240 (.Y(g8552),.A(g8217),.B(g8388));
OR2X1 OR2_241 (.Y(g5910),.A(g5023),.B(g4341));
OR2X1 OR2_242 (.Y(g11249),.A(g6162),.B(g11143));
OR2X1 OR2_243 (.Y(g11482),.A(g6628),.B(g11459));
OR2X1 OR_tmp232 (.Y(ttmp232),.A(g9410),.B(I14855));
OR2X1 OR_tmp233 (.Y(ttmp233),.A(g9612),.B(ttmp232));
OR2X1 OR_tmp234 (.Y(g9722),.A(g9643),.B(ttmp233));
OR2X1 OR_tmp235 (.Y(ttmp235),.A(g9933),.B(g9829));
OR2X1 OR_tmp236 (.Y(ttmp236),.A(g8168),.B(ttmp235));
OR2X1 OR_tmp237 (.Y(I15204),.A(g9904),.B(ttmp236));
OR2X1 OR2_244 (.Y(g7236),.A(g6684),.B(g6092));
OR2X1 OR_tmp238 (.Y(ttmp238),.A(g9205),.B(g9192));
OR2X1 OR_tmp239 (.Y(I14596),.A(g8995),.B(ttmp238));
OR2X1 OR2_245 (.Y(g8645),.A(g8127),.B(g8469));
OR2X1 OR2_246 (.Y(g11647),.A(g6622),.B(g11637));
OR2X1 OR2_247 (.Y(g6777),.A(g5691),.B(g5052));
OR2X1 OR_tmp240 (.Y(ttmp240),.A(g9658),.B(g9655));
OR2X1 OR_tmp241 (.Y(g9737),.A(g9657),.B(ttmp240));
OR2X1 OR_tmp242 (.Y(ttmp242),.A(g10468),.B(g10467));
OR2X1 OR_tmp243 (.Y(ttmp243),.A(g10472),.B(ttmp242));
OR2X1 OR_tmp244 (.Y(I16149),.A(g10470),.B(ttmp243));
OR2X1 OR2_248 (.Y(g11233),.A(g11085),.B(g10946));
OR2X1 OR2_249 (.Y(g8607),.A(g8406),.B(g8554));
OR2X1 OR_tmp245 (.Y(ttmp245),.A(g10476),.B(g10474));
OR2X1 OR_tmp246 (.Y(ttmp246),.A(g10386),.B(ttmp245));
OR2X1 OR_tmp247 (.Y(I16148),.A(g10384),.B(ttmp246));
OR2X1 OR2_250 (.Y(g8158),.A(g7893),.B(g6883));
OR2X1 OR2_251 (.Y(g5846),.A(g4932),.B(g4236));
OR2X1 OR2_252 (.Y(g5396),.A(g4481),.B(g3684));
OR2X1 OR2_253 (.Y(g5803),.A(g5575),.B(g4820));
OR2X1 OR2_254 (.Y(g11331),.A(g11272),.B(g11171));
OR2X1 OR2_255 (.Y(g7295),.A(g7071),.B(g6321));
OR2X1 OR2_256 (.Y(g6541),.A(g5788),.B(g5009));
OR2X1 OR2_257 (.Y(g8615),.A(g8413),.B(g8557));
OR2X1 OR2_258 (.Y(g9742),.A(g9173),.B(g9528));
OR2X1 OR2_259 (.Y(g9926),.A(g9868),.B(g9715));
OR2X1 OR2_260 (.Y(g9754),.A(g9173),.B(g9511));
OR2X1 OR2_261 (.Y(g8284),.A(g8102),.B(g7821));
OR2X1 OR2_262 (.Y(g2204),.A(g1393),.B(g1394));
OR2X1 OR2_263 (.Y(g7471),.A(g6880),.B(g6416));
OR2X1 OR2_264 (.Y(g7242),.A(g6693),.B(g6098));
OR2X1 OR2_265 (.Y(g5847),.A(g5626),.B(g4877));
OR2X1 OR2_266 (.Y(g6901),.A(g6788),.B(g6247));
OR2X1 OR2_267 (.Y(g8559),.A(g8380),.B(g4731));
OR2X1 OR_tmp248 (.Y(ttmp248),.A(g9357),.B(g9656));
OR2X1 OR_tmp249 (.Y(g9729),.A(g9618),.B(ttmp248));
OR2X1 OR2_268 (.Y(g10860),.A(g5513),.B(g10743));
OR2X1 OR2_269 (.Y(g9927),.A(g9869),.B(g9716));
OR2X1 OR2_270 (.Y(g10497),.A(g5052),.B(g10396));
OR2X1 OR_tmp250 (.Y(ttmp250),.A(g9662),.B(g9746));
OR2X1 OR_tmp251 (.Y(ttmp251),.A(g9739),.B(ttmp250));
OR2X1 OR_tmp252 (.Y(g9885),.A(g9598),.B(ttmp251));
OR2X1 OR_tmp253 (.Y(ttmp253),.A(g853),.B(g849));
OR2X1 OR_tmp254 (.Y(ttmp254),.A(g861),.B(ttmp253));
OR2X1 OR_tmp255 (.Y(g2528),.A(g857),.B(ttmp254));
OR2X1 OR2_271 (.Y(g11229),.A(g11154),.B(g11012));
OR2X1 OR2_272 (.Y(g8973),.A(g8821),.B(g8735));
OR2X1 OR2_273 (.Y(g10658),.A(g10595),.B(g7674));
OR2X1 OR2_274 (.Y(g10339),.A(g10232),.B(g9556));
OR2X1 OR_tmp256 (.Y(ttmp256),.A(g1157),.B(g1160));
OR2X1 OR_tmp257 (.Y(ttmp257),.A(g1149),.B(ttmp256));
OR2X1 OR_tmp258 (.Y(I5363),.A(g1153),.B(ttmp257));
OR2X1 OR2_275 (.Y(g11310),.A(g11220),.B(g11100));
OR2X1 OR2_276 (.Y(g6500),.A(g5725),.B(g4986));
OR2X1 OR2_277 (.Y(g10855),.A(g6075),.B(g10736));
OR2X1 OR2_278 (.Y(g9916),.A(g9855),.B(g9694));
OR2X1 OR2_279 (.Y(g10411),.A(g10299),.B(g9529));
OR2X1 OR2_280 (.Y(g11603),.A(g11582),.B(g11553));
OR2X1 OR_tmp259 (.Y(ttmp259),.A(g1255),.B(g1250));
OR2X1 OR_tmp260 (.Y(ttmp260),.A(g1265),.B(ttmp259));
OR2X1 OR_tmp261 (.Y(I5357),.A(g1260),.B(ttmp260));
OR2X1 OR2_281 (.Y(g9560),.A(g9052),.B(g9030));
OR2X1 OR2_282 (.Y(g6672),.A(g5941),.B(g5259));
OR2X1 OR_tmp262 (.Y(ttmp262),.A(g9599),.B(g9758));
OR2X1 OR_tmp263 (.Y(g9873),.A(g9623),.B(ttmp262));
OR2X1 OR2_283 (.Y(g6523),.A(g5745),.B(g4995));
OR2X1 OR2_284 (.Y(g10707),.A(g5545),.B(g10686));
OR2X1 OR_tmp264 (.Y(ttmp264),.A(g530),.B(g534));
OR2X1 OR_tmp265 (.Y(ttmp265),.A(g521),.B(ttmp264));
OR2X1 OR_tmp266 (.Y(I5626),.A(g525),.B(ttmp265));
OR2X1 OR2_285 (.Y(g9579),.A(g9052),.B(g9030));
OR2X1 OR2_286 (.Y(g7298),.A(g7136),.B(g6324));
OR2X1 OR2_287 (.Y(g6551),.A(g5804),.B(g5031));
OR2X1 OR2_288 (.Y(g6099),.A(g5273),.B(g4550));
OR2X1 OR2_289 (.Y(g8282),.A(g8101),.B(g7819));
OR2X1 OR2_290 (.Y(g9917),.A(g9856),.B(g9695));
OR2X1 OR_tmp267 (.Y(ttmp267),.A(g9624),.B(g9785));
OR2X1 OR_tmp268 (.Y(ttmp268),.A(g7853),.B(ttmp267));
OR2X1 OR_tmp269 (.Y(I15057),.A(g9680),.B(ttmp268));
OR2X1 OR2_291 (.Y(g7219),.A(g6661),.B(g6076));
OR2X1 OR2_292 (.Y(g10019),.A(I15219),.B(I15220));
OR2X1 OR2_293 (.Y(g5857),.A(g5418),.B(g4670));
OR2X1 OR_tmp270 (.Y(ttmp270),.A(g9616),.B(I14862));
OR2X1 OR_tmp271 (.Y(ttmp271),.A(g9642),.B(ttmp270));
OR2X1 OR_tmp272 (.Y(g9725),.A(g9659),.B(ttmp271));
OR2X1 OR2_294 (.Y(g11298),.A(g11212),.B(g11087));
OR2X1 OR2_295 (.Y(g10402),.A(g10295),.B(g9554));
OR2X1 OR_tmp273 (.Y(ttmp273),.A(g476),.B(I5626));
OR2X1 OR_tmp274 (.Y(ttmp274),.A(g538),.B(ttmp273));
OR2X1 OR_tmp275 (.Y(g2521),.A(g542),.B(ttmp274));
OR2X1 OR_tmp276 (.Y(ttmp276),.A(g9205),.B(g9192));
OR2X1 OR_tmp277 (.Y(I14751),.A(g8995),.B(ttmp276));
OR2X1 OR2_296 (.Y(g10866),.A(g5539),.B(g10753));
OR2X1 OR2_297 (.Y(g6534),.A(g5772),.B(g5003));
OR2X1 OR2_298 (.Y(g11232),.A(g11158),.B(g11015));
OR2X1 OR_tmp278 (.Y(ttmp278),.A(g9386),.B(g9591));
OR2X1 OR_tmp279 (.Y(g9706),.A(g9644),.B(ttmp278));
OR2X1 OR2_299 (.Y(g10001),.A(I15204),.B(I15205));
OR2X1 OR2_300 (.Y(g8776),.A(g5510),.B(g8655));
OR2X1 OR2_301 (.Y(g7225),.A(g6666),.B(g6079));
OR2X1 OR_tmp280 (.Y(ttmp280),.A(g9608),.B(g9757));
OR2X1 OR_tmp281 (.Y(g9888),.A(g9648),.B(ttmp280));
OR2X1 OR2_302 (.Y(g11261),.A(g11238),.B(g11023));
OR2X1 OR_tmp282 (.Y(ttmp282),.A(g9942),.B(g9815));
OR2X1 OR_tmp283 (.Y(g9956),.A(g9948),.B(ttmp282));
OR2X1 OR2_303 (.Y(g10923),.A(g10778),.B(g10715));
OR2X1 OR2_304 (.Y(g8264),.A(g7879),.B(g3389));
OR2X1 OR2_305 (.Y(g6513),.A(g5737),.B(g4991));
OR2X1 OR_tmp284 (.Y(ttmp284),.A(g9645),.B(g9588));
OR2X1 OR_tmp285 (.Y(I14835),.A(g9621),.B(ttmp284));
OR2X1 OR2_306 (.Y(g8641),.A(g8120),.B(g8463));
OR2X1 OR_tmp286 (.Y(ttmp286),.A(g4093),.B(g126));
OR2X1 OR_tmp287 (.Y(g5361),.A(g4316),.B(ttmp286));
OR2X1 OR2_307 (.Y(g11316),.A(g11226),.B(g11103));
OR2X1 OR_tmp288 (.Y(ttmp288),.A(g10477),.B(g10475));
OR2X1 OR_tmp289 (.Y(ttmp289),.A(g10479),.B(ttmp288));
OR2X1 OR_tmp290 (.Y(I16161),.A(g10478),.B(ttmp289));
OR2X1 OR2_308 (.Y(g6916),.A(g6348),.B(g5687));
OR2X1 OR2_309 (.Y(g8777),.A(g5522),.B(g8659));
OR2X1 OR_tmp291 (.Y(ttmp291),.A(g1411),.B(g1415));
OR2X1 OR_tmp292 (.Y(ttmp292),.A(g1403),.B(ttmp291));
OR2X1 OR_tmp293 (.Y(g2353),.A(g1407),.B(ttmp292));
OR2X1 OR2_310 (.Y(g7510),.A(g7186),.B(g6730));
OR2X1 OR_tmp294 (.Y(ttmp294),.A(g9943),.B(g9776));
OR2X1 OR_tmp295 (.Y(g9957),.A(g9949),.B(ttmp294));
OR2X1 OR2_311 (.Y(g2744),.A(I5804),.B(I5805));
OR2X1 OR2_312 (.Y(g7245),.A(g6696),.B(g6102));
OR2X1 OR2_313 (.Y(g7291),.A(g7050),.B(g6317));
OR2X1 OR2_314 (.Y(g8611),.A(g8410),.B(g8556));
OR2X1 OR_tmp296 (.Y(ttmp296),.A(g9932),.B(g9828));
OR2X1 OR_tmp297 (.Y(ttmp297),.A(g8167),.B(ttmp296));
OR2X1 OR_tmp298 (.Y(I15199),.A(g9903),.B(ttmp297));
OR2X1 OR2_315 (.Y(g10550),.A(g4942),.B(g10450));
OR2X1 OR2_316 (.Y(g11330),.A(g11304),.B(g11170));
OR2X1 OR2_317 (.Y(g10721),.A(g10306),.B(g10669));
OR2X1 OR2_318 (.Y(g8153),.A(g7888),.B(g6875));
OR2X1 OR2_319 (.Y(g10773),.A(g5540),.B(g10685));
OR2X1 OR2_320 (.Y(g3688),.A(g3144),.B(g2454));
OR2X1 OR_tmp299 (.Y(ttmp299),.A(g9859),.B(g9881));
OR2X1 OR_tmp300 (.Y(ttmp300),.A(g9842),.B(ttmp299));
OR2X1 OR_tmp301 (.Y(I15225),.A(g9967),.B(ttmp300));
OR2X1 OR2_321 (.Y(g6042),.A(g5535),.B(g3987));
OR2X1 OR2_322 (.Y(g10655),.A(g10561),.B(g7389));
OR2X1 OR2_323 (.Y(g11259),.A(g11236),.B(g11021));
OR2X1 OR2_324 (.Y(g11225),.A(g11149),.B(g11009));
OR2X1 OR2_325 (.Y(g5914),.A(g5029),.B(g4343));
OR2X1 OR2_326 (.Y(g11258),.A(g11235),.B(g11020));
OR2X1 OR2_327 (.Y(g6054),.A(g5199),.B(g4483));
OR2X1 OR_tmp302 (.Y(ttmp302),.A(g9422),.B(g9426));
OR2X1 OR_tmp303 (.Y(g9728),.A(g9412),.B(ttmp302));
OR2X1 OR_tmp304 (.Y(ttmp304),.A(g9425),.B(g9423));
OR2X1 OR_tmp305 (.Y(g9730),.A(g9414),.B(ttmp304));
OR2X1 OR2_328 (.Y(g5820),.A(g5595),.B(g4834));
OR2X1 OR_tmp306 (.Y(ttmp306),.A(g7853),.B(g8465));
OR2X1 OR_tmp307 (.Y(g8574),.A(g5679),.B(ttmp306));
OR2X1 OR2_329 (.Y(g11602),.A(g11581),.B(g11552));
OR2X1 OR2_330 (.Y(g10502),.A(g4169),.B(g10365));
OR2X1 OR2_331 (.Y(g10557),.A(g4123),.B(g10508));
OR2X1 OR_tmp308 (.Y(ttmp308),.A(g9896),.B(g9835));
OR2X1 OR_tmp309 (.Y(ttmp309),.A(g8175),.B(ttmp308));
OR2X1 OR_tmp310 (.Y(I15171),.A(g9909),.B(ttmp309));
OR2X1 OR2_332 (.Y(g11337),.A(g11282),.B(g11177));
OR2X1 OR2_333 (.Y(g7465),.A(g6876),.B(g6410));
OR2X1 OR2_334 (.Y(g8262),.A(g7970),.B(g7625));
OR2X1 OR2_335 (.Y(g8889),.A(g8844),.B(g8756));
OR2X1 OR2_336 (.Y(g7096),.A(g6544),.B(g5911));
OR2X1 OR2_337 (.Y(g5995),.A(g5097),.B(g5099));
OR2X1 OR2_338 (.Y(g8285),.A(g8104),.B(g7822));
OR2X1 OR2_339 (.Y(g10791),.A(g6186),.B(g10762));
OR2X1 OR2_340 (.Y(g2499),.A(I5570),.B(I5571));
OR2X1 OR_tmp311 (.Y(ttmp311),.A(g9205),.B(g9192));
OR2X1 OR_tmp312 (.Y(I14607),.A(g8995),.B(ttmp311));
OR2X1 OR2_341 (.Y(g6049),.A(g5254),.B(g3718));
OR2X1 OR2_342 (.Y(g9920),.A(g9860),.B(g9701));
OR2X1 OR2_343 (.Y(g10556),.A(g4115),.B(g10506));
OR2X1 OR2_344 (.Y(g8643),.A(g8364),.B(g8508));
OR2X1 OR2_345 (.Y(g5810),.A(g5588),.B(g4823));
OR2X1 OR2_346 (.Y(g11336),.A(g11281),.B(g11176));
OR2X1 OR2_347 (.Y(g8742),.A(g8135),.B(g8598));
OR2X1 OR2_348 (.Y(g8926),.A(g8848),.B(g8764));
OR2X1 OR2_349 (.Y(g7218),.A(g6655),.B(g6070));
OR2X1 OR_tmp313 (.Y(ttmp313),.A(g9937),.B(g9834));
OR2X1 OR_tmp314 (.Y(ttmp314),.A(g8174),.B(ttmp313));
OR2X1 OR_tmp315 (.Y(I15224),.A(g9908),.B(ttmp314));
OR2X1 OR2_350 (.Y(g7293),.A(g7063),.B(g6319));
OR2X1 OR2_351 (.Y(g11288),.A(g11204),.B(g11070));
OR2X1 OR2_352 (.Y(g10800),.A(g6245),.B(g10772));
OR2X1 OR2_353 (.Y(g11308),.A(g11218),.B(g11098));
OR2X1 OR2_354 (.Y(g8269),.A(g7892),.B(g3429));
OR2X1 OR2_355 (.Y(g10417),.A(g10301),.B(g9527));
OR2X1 OR2_356 (.Y(g10936),.A(g5170),.B(g10808));
OR2X1 OR2_357 (.Y(g9388),.A(g9240),.B(g9223));
OR2X1 OR2_358 (.Y(g6185),.A(g5470),.B(g4715));
OR2X1 OR2_359 (.Y(g6470),.A(g5699),.B(g4960));
OR2X1 OR2_360 (.Y(g6897),.A(g6771),.B(g6240));
OR2X1 OR2_361 (.Y(g8885),.A(g8841),.B(g8754));
OR2X1 OR2_362 (.Y(g11260),.A(g11237),.B(g11022));
OR2X1 OR2_363 (.Y(g11488),.A(g6671),.B(g11465));
OR2X1 OR2_364 (.Y(g6105),.A(g5279),.B(g4559));
OR2X1 OR2_365 (.Y(g10807),.A(g10701),.B(g10761));
OR2X1 OR2_366 (.Y(g10639),.A(g10623),.B(g7734));
OR2X1 OR2_367 (.Y(g4556),.A(g3536),.B(g2916));
OR2X1 OR2_368 (.Y(g8288),.A(g8119),.B(g7825));
OR2X1 OR2_369 (.Y(g6755),.A(g6106),.B(g5479));
OR2X1 OR_tmp316 (.Y(ttmp316),.A(g9600),.B(g9611));
OR2X1 OR_tmp317 (.Y(I14862),.A(g9587),.B(ttmp316));
OR2X1 OR_tmp318 (.Y(ttmp318),.A(g10482),.B(g10481));
OR2X1 OR_tmp319 (.Y(ttmp319),.A(g10394),.B(ttmp318));
OR2X1 OR_tmp320 (.Y(I16160),.A(g10392),.B(ttmp319));
OR2X1 OR_tmp321 (.Y(ttmp321),.A(g9624),.B(g9785));
OR2X1 OR_tmp322 (.Y(ttmp322),.A(g7853),.B(ttmp321));
OR2X1 OR_tmp323 (.Y(I15042),.A(g9686),.B(ttmp322));
OR2X1 OR2_370 (.Y(g11610),.A(g11589),.B(g11560));
OR2X1 OR_tmp324 (.Y(ttmp324),.A(g9359),.B(g9589));
OR2X1 OR_tmp325 (.Y(ttmp325),.A(g9660),.B(ttmp324));
OR2X1 OR_tmp326 (.Y(g9711),.A(g9390),.B(ttmp325));
OR2X1 OR2_371 (.Y(g6045),.A(g5541),.B(g3989));
OR2X1 OR2_372 (.Y(g11270),.A(g11198),.B(g11032));
OR2X1 OR2_373 (.Y(g7258),.A(g6549),.B(g5913));
OR2X1 OR2_374 (.Y(g6059),.A(g5211),.B(g4489));
OR2X1 OR2_375 (.Y(g10007),.A(I15209),.B(I15210));
OR2X1 OR2_376 (.Y(g11267),.A(g11192),.B(g11029));
OR2X1 OR2_377 (.Y(g11294),.A(g6576),.B(g11210));
OR2X1 OR_tmp327 (.Y(ttmp327),.A(g9125),.B(g9111));
OR2X1 OR_tmp328 (.Y(g9509),.A(g9151),.B(ttmp327));
OR2X1 OR2_378 (.Y(g7211),.A(g6647),.B(g6067));
OR2X1 OR2_379 (.Y(g5404),.A(g4487),.B(g3696));
OR2X1 OR2_380 (.Y(g4089),.A(g1959),.B(g3318));
OR2X1 OR_tmp329 (.Y(ttmp329),.A(g9936),.B(g9833));
OR2X1 OR_tmp330 (.Y(ttmp330),.A(g8172),.B(ttmp329));
OR2X1 OR_tmp331 (.Y(I15219),.A(g9907),.B(ttmp330));
OR2X1 OR2_381 (.Y(g11219),.A(g11145),.B(g11006));
OR2X1 OR2_382 (.Y(g6015),.A(g5497),.B(g3942));
OR2X1 OR2_383 (.Y(g10720),.A(g10304),.B(g10667));
OR2X1 OR2_384 (.Y(g8265),.A(g7881),.B(g3396));
OR2X1 OR2_385 (.Y(g5224),.A(g4360),.B(g3512));
OR2X1 OR_tmp332 (.Y(ttmp332),.A(g9667),.B(I14827));
OR2X1 OR_tmp333 (.Y(g9700),.A(g9358),.B(ttmp332));
OR2X1 OR2_386 (.Y(g7106),.A(g6554),.B(g5917));
OR2X1 OR2_387 (.Y(g8770),.A(g5476),.B(g8651));
OR2X1 OR2_388 (.Y(g11201),.A(g11152),.B(g11011));
OR2X1 OR_tmp334 (.Y(ttmp334),.A(g9898),.B(g9779));
OR2X1 OR_tmp335 (.Y(g9950),.A(g9901),.B(ttmp334));
OR2X1 OR_tmp336 (.Y(ttmp336),.A(g9391),.B(I14858));
OR2X1 OR_tmp337 (.Y(ttmp337),.A(g9620),.B(ttmp336));
OR2X1 OR_tmp338 (.Y(g9723),.A(g9652),.B(ttmp337));
OR2X1 OR2_389 (.Y(g2309),.A(I5357),.B(I5358));
OR2X1 OR2_390 (.Y(g11266),.A(g11190),.B(g11028));
OR2X1 OR2_391 (.Y(g10727),.A(g4969),.B(g10638));
OR2X1 OR2_392 (.Y(g10863),.A(g5531),.B(g10750));
OR2X1 OR2_393 (.Y(g8429),.A(g8385),.B(g8069));
OR2X1 OR2_394 (.Y(g9751),.A(g9515),.B(g9510));
OR2X1 OR2_395 (.Y(g8281),.A(g8097),.B(g7818));
OR2X1 OR2_396 (.Y(g6910),.A(g6341),.B(g5680));
OR2X1 OR2_397 (.Y(g8639),.A(g8118),.B(g8462));
OR2X1 OR_tmp339 (.Y(ttmp339),.A(g9292),.B(g9274));
OR2X1 OR_tmp340 (.Y(g9673),.A(g9454),.B(ttmp339));
OR2X1 OR2_398 (.Y(g11285),.A(g11255),.B(g11161));
OR2X1 OR2_399 (.Y(g11305),.A(g11215),.B(g11093));
OR2X1 OR_tmp341 (.Y(ttmp341),.A(g9863),.B(g9876));
OR2X1 OR_tmp342 (.Y(ttmp342),.A(g9844),.B(ttmp341));
OR2X1 OR_tmp343 (.Y(I15177),.A(g9960),.B(ttmp342));
OR2X1 OR_tmp344 (.Y(ttmp344),.A(g9428),.B(g9421));
OR2X1 OR_tmp345 (.Y(g9734),.A(g9415),.B(ttmp344));
OR2X1 OR_tmp346 (.Y(ttmp346),.A(g9614),.B(g9584));
OR2X1 OR_tmp347 (.Y(I14827),.A(g9603),.B(ttmp346));
OR2X1 OR2_400 (.Y(g5824),.A(g5602),.B(g4839));
OR2X1 OR2_401 (.Y(g8715),.A(g8416),.B(g8687));
OR2X1 OR2_402 (.Y(g5762),.A(g5178),.B(g5186));
OR2X1 OR2_403 (.Y(g6538),.A(g5782),.B(g5006));
OR2X1 OR2_404 (.Y(g5590),.A(g4718),.B(g4723));
OR2X1 OR2_405 (.Y(g10726),.A(g10316),.B(g10673));
OR2X1 OR2_406 (.Y(g3120),.A(I6350),.B(I6351));
OR2X1 OR2_407 (.Y(g9573),.A(g9052),.B(g9030));
OR2X1 OR_tmp348 (.Y(ttmp348),.A(g3563),.B(g1527));
OR2X1 OR_tmp349 (.Y(g4640),.A(g3348),.B(ttmp348));
OR2X1 OR2_408 (.Y(g6093),.A(g5264),.B(g4534));
OR2X1 OR2_409 (.Y(g8162),.A(g7898),.B(g6889));
OR2X1 OR2_410 (.Y(g8268),.A(g7962),.B(g7613));
OR2X1 OR2_411 (.Y(g9569),.A(g9052),.B(g9030));
OR2X1 OR2_412 (.Y(g11485),.A(g6646),.B(g11462));
OR2X1 OR2_413 (.Y(g10797),.A(g6206),.B(g10766));
OR2X1 OR_tmp350 (.Y(ttmp350),.A(g9205),.B(g9192));
OR2X1 OR_tmp351 (.Y(I14779),.A(g8995),.B(ttmp350));
OR2X1 OR2_414 (.Y(g10408),.A(g10298),.B(g9553));
OR2X1 OR2_415 (.Y(g10635),.A(g10622),.B(g7732));
OR2X1 OR2_416 (.Y(g2305),.A(I5351),.B(I5352));
OR2X1 OR_tmp352 (.Y(ttmp352),.A(g9897),.B(g9836));
OR2X1 OR_tmp353 (.Y(ttmp353),.A(g8176),.B(ttmp352));
OR2X1 OR_tmp354 (.Y(I15176),.A(g9910),.B(ttmp353));
OR2X1 OR2_417 (.Y(g3435),.A(g2945),.B(g2950));
OR2X1 OR2_418 (.Y(g9924),.A(g9866),.B(g9709));
OR2X1 OR2_419 (.Y(g10711),.A(g5547),.B(g10690));
OR2X1 OR2_420 (.Y(g5814),.A(g5591),.B(g4827));
OR2X1 OR2_421 (.Y(g5038),.A(g4878),.B(g4884));
OR2X1 OR_tmp355 (.Y(ttmp355),.A(g9854),.B(g9879));
OR2X1 OR_tmp356 (.Y(ttmp356),.A(g9840),.B(ttmp355));
OR2X1 OR_tmp357 (.Y(I15215),.A(g9965),.B(ttmp356));
OR2X1 OR2_422 (.Y(g8226),.A(g7504),.B(g8002));
OR2X1 OR2_423 (.Y(g7367),.A(g7224),.B(g6744));
OR2X1 OR2_424 (.Y(g7457),.A(g6873),.B(g6404));
OR2X1 OR2_425 (.Y(g5229),.A(g4364),.B(g3516));
OR2X1 OR2_426 (.Y(g5993),.A(g5090),.B(g4400));
OR2X1 OR2_427 (.Y(g8283),.A(g8098),.B(g7820));
OR2X1 OR2_428 (.Y(g7971),.A(g5110),.B(g7549));
OR2X1 OR2_429 (.Y(g8602),.A(g8401),.B(g8550));
OR2X1 OR2_430 (.Y(g8920),.A(g8845),.B(g8759));
OR2X1 OR2_431 (.Y(g10663),.A(g10237),.B(g10581));
OR2X1 OR2_432 (.Y(g6074),.A(g5349),.B(g1));
OR2X1 OR2_433 (.Y(g8261),.A(g7876),.B(g3383));
OR2X1 OR2_434 (.Y(g10862),.A(g5524),.B(g10746));
OR2X1 OR2_435 (.Y(g5837),.A(g5640),.B(g4224));
OR2X1 OR2_436 (.Y(g11333),.A(g11274),.B(g11173));
OR2X1 OR2_437 (.Y(g6080),.A(g5249),.B(g4512));
OR2X1 OR2_438 (.Y(g6480),.A(g5721),.B(g4971));
OR2X1 OR2_439 (.Y(g7740),.A(g7209),.B(g6741));
OR2X1 OR2_440 (.Y(g10702),.A(g10562),.B(g3877));
OR2X1 OR_tmp358 (.Y(ttmp358),.A(g9606),.B(I14822));
OR2X1 OR_tmp359 (.Y(g9697),.A(g9665),.B(ttmp358));
OR2X1 OR2_441 (.Y(g8203),.A(g7453),.B(g7999));
OR2X1 OR2_442 (.Y(g9914),.A(g9851),.B(g9692));
OR2X1 OR2_443 (.Y(g10564),.A(g10560),.B(g7368));
OR2X1 OR2_444 (.Y(g11484),.A(g6639),.B(g11461));
OR2X1 OR2_445 (.Y(g5842),.A(g5618),.B(g4870));
OR2X1 OR_tmp360 (.Y(ttmp360),.A(g9848),.B(g9880));
OR2X1 OR_tmp361 (.Y(ttmp361),.A(g9837),.B(ttmp360));
OR2X1 OR_tmp362 (.Y(I15200),.A(g9962),.B(ttmp361));
OR2X1 OR2_446 (.Y(g11609),.A(g11588),.B(g11559));
OR2X1 OR_tmp363 (.Y(ttmp363),.A(g9205),.B(g9192));
OR2X1 OR_tmp364 (.Y(I14582),.A(g8995),.B(ttmp363));
OR2X1 OR2_447 (.Y(g8940),.A(g8793),.B(g8703));
OR2X1 OR2_448 (.Y(g11312),.A(g11222),.B(g11101));
OR2X1 OR2_449 (.Y(g11608),.A(g11587),.B(g11558));
OR2X1 OR2_450 (.Y(g6000),.A(g5480),.B(g3912));
OR2X1 OR2_451 (.Y(g8428),.A(g8382),.B(g8068));
OR2X1 OR2_452 (.Y(g8430),.A(g8386),.B(g8070));
OR2X1 OR2_453 (.Y(g9922),.A(g9864),.B(g9705));
OR2X1 OR2_454 (.Y(g8247),.A(g8010),.B(g7704));
OR2X1 OR2_455 (.Y(g3438),.A(g2939),.B(g2944));
OR2X1 OR_tmp365 (.Y(ttmp365),.A(g440),.B(g444));
OR2X1 OR_tmp366 (.Y(ttmp366),.A(g431),.B(ttmp365));
OR2X1 OR_tmp367 (.Y(I5576),.A(g435),.B(ttmp366));
OR2X1 OR2_456 (.Y(g6924),.A(g6362),.B(g4261));
OR2X1 OR2_457 (.Y(g5405),.A(g4476),.B(g3440));
OR2X1 OR2_458 (.Y(g8638),.A(g8108),.B(g8461));
OR2X1 OR2_459 (.Y(g8609),.A(g8408),.B(g8555));
OR2X1 OR2_460 (.Y(g9995),.A(I15199),.B(I15200));
OR2X1 OR2_461 (.Y(g8883),.A(g8838),.B(g8753));
OR2X1 OR_tmp368 (.Y(ttmp368),.A(g9935),.B(g9831));
OR2X1 OR_tmp369 (.Y(ttmp369),.A(g8170),.B(ttmp368));
OR2X1 OR_tmp370 (.Y(I15214),.A(g9906),.B(ttmp369));
OR2X1 OR_tmp371 (.Y(ttmp371),.A(g1458),.B(I5649));
OR2X1 OR_tmp372 (.Y(g2538),.A(g1466),.B(ttmp371));
OR2X1 OR2_462 (.Y(g11329),.A(g11302),.B(g11169));
OR2X1 OR2_463 (.Y(g4255),.A(g4009),.B(g4047));
OR2X1 OR2_464 (.Y(g11328),.A(g11299),.B(g11168));
OR2X1 OR_tmp373 (.Y(ttmp373),.A(g9605),.B(I14835));
OR2X1 OR_tmp374 (.Y(g9704),.A(g9385),.B(ttmp373));
OR2X1 OR_tmp375 (.Y(ttmp375),.A(g1121),.B(g1117));
OR2X1 OR_tmp376 (.Y(ttmp376),.A(g1129),.B(ttmp375));
OR2X1 OR_tmp377 (.Y(I5352),.A(g1125),.B(ttmp376));
OR2X1 OR2_465 (.Y(g8774),.A(g5499),.B(g8654));
OR2X1 OR_tmp378 (.Y(ttmp378),.A(g9940),.B(g9781));
OR2X1 OR_tmp379 (.Y(g9954),.A(g9946),.B(ttmp378));
OR2X1 OR2_466 (.Y(g10405),.A(g10297),.B(g9530));
OR2X1 OR2_467 (.Y(g9363),.A(g9205),.B(g9192));
OR2X1 OR2_468 (.Y(g5849),.A(g4949),.B(g4260));
OR2X1 OR_tmp380 (.Y(ttmp380),.A(g506),.B(g501));
OR2X1 OR_tmp381 (.Y(ttmp381),.A(g516),.B(ttmp380));
OR2X1 OR_tmp382 (.Y(I5599),.A(g511),.B(ttmp381));
OR2X1 OR2_469 (.Y(g7204),.A(g6645),.B(g6062));
OR2X1 OR2_470 (.Y(g7300),.A(g7139),.B(g6326));
OR2X1 OR2_471 (.Y(g4293),.A(g4064),.B(g4068));
OR2X1 OR2_472 (.Y(g9912),.A(g9847),.B(g9690));
OR2X1 OR2_473 (.Y(g6533),.A(g5771),.B(g5002));
OR2X1 OR2_474 (.Y(g8816),.A(g7951),.B(g8731));
OR2X1 OR2_475 (.Y(g9929),.A(g9871),.B(g9718));
OR2X1 OR2_476 (.Y(g5819),.A(g5625),.B(g4876));
OR2X1 OR_tmp383 (.Y(ttmp383),.A(g9622),.B(g9586));
OR2X1 OR_tmp384 (.Y(I14831),.A(g9613),.B(ttmp383));
OR2X1 OR2_477 (.Y(g5852),.A(g5632),.B(g4883));
OR2X1 OR2_478 (.Y(g8263),.A(g8032),.B(g7720));
OR2X1 OR2_479 (.Y(g3431),.A(g2951),.B(g2957));
OR2X1 OR_tmp385 (.Y(ttmp385),.A(g9292),.B(g9274));
OR2X1 OR_tmp386 (.Y(g9683),.A(g9454),.B(ttmp385));
OR2X1 OR2_480 (.Y(g8631),.A(g8474),.B(g7449));
OR2X1 OR2_481 (.Y(g6922),.A(g6352),.B(g5694));
OR2X1 OR2_482 (.Y(g8817),.A(g7954),.B(g8732));
OR2X1 OR_tmp387 (.Y(ttmp387),.A(g9384),.B(g9361));
OR2X1 OR_tmp388 (.Y(ttmp388),.A(g9649),.B(ttmp387));
OR2X1 OR_tmp389 (.Y(g9735),.A(g9651),.B(ttmp388));
OR2X1 OR2_483 (.Y(g8605),.A(g8404),.B(g8553));
OR2X1 OR2_484 (.Y(g11263),.A(g11187),.B(g11025));
OR2X1 OR2_485 (.Y(g6739),.A(g5769),.B(g5780));
OR2X1 OR2_486 (.Y(g11332),.A(g11273),.B(g11172));
OR2X1 OR2_487 (.Y(g7143),.A(g6619),.B(g6039));
OR2X1 OR2_488 (.Y(g6479),.A(g5707),.B(g4968));
OR2X1 OR_tmp390 (.Y(ttmp390),.A(g9624),.B(g9785));
OR2X1 OR_tmp391 (.Y(ttmp391),.A(g7853),.B(ttmp390));
OR2X1 OR_tmp392 (.Y(I15048),.A(g9683),.B(ttmp391));
OR2X1 OR2_489 (.Y(g6501),.A(g5726),.B(g4987));
OR2X1 OR_tmp393 (.Y(ttmp393),.A(g9647),.B(I14831));
OR2X1 OR_tmp394 (.Y(g9702),.A(g9365),.B(ttmp393));
OR2X1 OR2_490 (.Y(g11221),.A(g11146),.B(g11007));
OR2X1 OR_tmp395 (.Y(ttmp395),.A(g9938),.B(g9817));
OR2X1 OR_tmp396 (.Y(g9952),.A(g9944),.B(ttmp395));
OR2X1 OR2_491 (.Y(g11613),.A(g11600),.B(g11591));
OR2X1 OR2_492 (.Y(g7621),.A(g5108),.B(g6994));
OR2X1 OR2_493 (.Y(g3399),.A(g2918),.B(g2940));
OR2X1 OR2_494 (.Y(g11605),.A(g11584),.B(g11555));
OR2X1 OR2_495 (.Y(g4274),.A(g4054),.B(g4058));
OR2X1 OR_tmp397 (.Y(ttmp397),.A(g9205),.B(g9192));
OR2X1 OR_tmp398 (.Y(I14602),.A(g8995),.B(ttmp397));
OR2X1 OR_tmp399 (.Y(ttmp399),.A(g9624),.B(g9785));
OR2X1 OR_tmp400 (.Y(ttmp400),.A(g7853),.B(ttmp399));
OR2X1 OR_tmp401 (.Y(I15033),.A(g9804),.B(ttmp400));
OR2X1 OR2_496 (.Y(g10717),.A(g6235),.B(g10705));
OR2X1 OR_tmp402 (.Y(ttmp402),.A(g841),.B(g837));
OR2X1 OR_tmp403 (.Y(I5629),.A(g845),.B(ttmp402));
OR2X1 OR2_497 (.Y(g9925),.A(g9867),.B(g9712));
OR2X1 OR2_498 (.Y(g3819),.A(g3275),.B(g9));
OR2X1 OR2_499 (.Y(g6912),.A(g6350),.B(g4235));
OR2X1 OR2_500 (.Y(g10723),.A(g4952),.B(g10633));
OR2X1 OR2_501 (.Y(g6929),.A(g6360),.B(g5704));
OR2X1 OR2_502 (.Y(g10646),.A(g10625),.B(g7739));
OR2X1 OR2_503 (.Y(g9516),.A(g9151),.B(g9125));
OR2X1 OR2_504 (.Y(g6626),.A(g5934),.B(g123));
OR2X1 OR_tmp404 (.Y(ttmp404),.A(g2433),.B(g2419));
OR2X1 OR_tmp405 (.Y(ttmp405),.A(g2445),.B(ttmp404));
OR2X1 OR_tmp406 (.Y(I6350),.A(g2437),.B(ttmp405));
OR2X1 OR2_505 (.Y(g11325),.A(g11295),.B(g11165));
OR2X1 OR_tmp407 (.Y(ttmp407),.A(g1292),.B(g1296));
OR2X1 OR_tmp408 (.Y(ttmp408),.A(g1280),.B(ttmp407));
OR2X1 OR_tmp409 (.Y(I5366),.A(g1284),.B(ttmp408));
OR2X1 OR_tmp410 (.Y(ttmp410),.A(g1486),.B(g1482));
OR2X1 OR_tmp411 (.Y(I5649),.A(g1499),.B(ttmp410));
OR2X1 OR2_506 (.Y(g6894),.A(g6763),.B(g4868));
OR2X1 OR_tmp412 (.Y(ttmp412),.A(g9447),.B(g9506));
OR2X1 OR_tmp413 (.Y(g9738),.A(g9417),.B(ttmp412));
OR2X1 OR2_507 (.Y(g8383),.A(g8163),.B(g5051));
OR2X1 OR2_508 (.Y(g8779),.A(g5530),.B(g8663));
OR2X1 OR2_509 (.Y(g8161),.A(g8005),.B(g7185));
OR2X1 OR2_510 (.Y(g8451),.A(g3440),.B(g8366));
OR2X1 OR2_511 (.Y(g9915),.A(g9853),.B(g9693));
OR2X1 OR_tmp414 (.Y(ttmp414),.A(g1270),.B(I5366));
OR2X1 OR_tmp415 (.Y(ttmp415),.A(g1300),.B(ttmp414));
OR2X1 OR_tmp416 (.Y(g2316),.A(g1304),.B(ttmp415));
OR2X1 OR2_512 (.Y(g5576),.A(g4675),.B(g3664));
OR2X1 OR2_513 (.Y(g10857),.A(g6090),.B(g10738));
OR2X1 OR2_514 (.Y(g10793),.A(g6194),.B(g10763));
OR2X1 OR2_515 (.Y(g7511),.A(g6890),.B(g6438));
OR2X1 OR2_516 (.Y(g8944),.A(g8799),.B(g8708));
OR2X1 OR2_517 (.Y(g10765),.A(g5492),.B(g10680));
OR2X1 OR2_518 (.Y(g10549),.A(g4951),.B(g10451));
OR2X1 OR2_519 (.Y(g7092),.A(g6540),.B(g5902));
OR2X1 OR2_520 (.Y(g11604),.A(g11583),.B(g11554));
OR2X1 OR2_521 (.Y(g8434),.A(g8400),.B(g8074));
OR2X1 OR2_522 (.Y(g6546),.A(g5796),.B(g5026));
OR2X1 OR2_523 (.Y(g3354),.A(g2920),.B(g2124));
OR2X1 OR2_524 (.Y(g9928),.A(g9870),.B(g9717));
OR2X1 OR2_525 (.Y(g11262),.A(g11240),.B(g11024));
OR2X1 OR_tmp417 (.Y(ttmp417),.A(g9388),.B(g9363));
OR2X1 OR_tmp418 (.Y(ttmp418),.A(g9010),.B(ttmp417));
OR2X1 OR_tmp419 (.Y(g9785),.A(g8995),.B(ttmp418));
OR2X1 OR2_526 (.Y(g5867),.A(g3440),.B(g4921));
OR2X1 OR2_527 (.Y(g8210),.A(g7466),.B(g7995));
OR2X1 OR2_528 (.Y(g10533),.A(g4933),.B(g10449));
OR2X1 OR2_529 (.Y(g9563),.A(g9052),.B(g9030));
OR2X1 OR2_530 (.Y(g6906),.A(g6791),.B(g5674));
OR2X1 OR2_531 (.Y(g7375),.A(g7230),.B(g6745));
OR2X1 OR2_532 (.Y(g7651),.A(g7135),.B(g4084));
OR2X1 OR_tmp420 (.Y(ttmp420),.A(g406),.B(g401));
OR2X1 OR_tmp421 (.Y(ttmp421),.A(g416),.B(ttmp420));
OR2X1 OR_tmp422 (.Y(I5570),.A(g411),.B(ttmp421));
OR2X1 OR_tmp423 (.Y(ttmp423),.A(g9364),.B(g9387));
OR2X1 OR_tmp424 (.Y(g9731),.A(g9641),.B(ttmp423));
OR2X1 OR2_533 (.Y(g11247),.A(g11097),.B(g10949));
OR2X1 OR_tmp425 (.Y(ttmp425),.A(g9624),.B(g9785));
OR2X1 OR_tmp426 (.Y(ttmp426),.A(g7853),.B(ttmp425));
OR2X1 OR_tmp427 (.Y(I15045),.A(g9676),.B(ttmp426));
OR2X1 OR2_534 (.Y(g10856),.A(g6083),.B(g10737));
OR2X1 OR2_535 (.Y(g9557),.A(g9052),.B(g9030));
OR2X1 OR2_536 (.Y(g7184),.A(g6625),.B(g6047));
OR2X1 OR2_537 (.Y(g11612),.A(g11599),.B(g11590));
OR2X1 OR2_538 (.Y(g7384),.A(g7088),.B(g6618));
OR2X1 OR2_539 (.Y(g11324),.A(g11271),.B(g11164));
OR2X1 OR2_540 (.Y(g8922),.A(g8822),.B(g8736));
OR2X1 OR_tmp428 (.Y(ttmp428),.A(g1235),.B(g1275));
OR2X1 OR_tmp429 (.Y(ttmp429),.A(g1245),.B(ttmp428));
OR2X1 OR_tmp430 (.Y(I5358),.A(g1240),.B(ttmp429));
OR2X1 OR_tmp431 (.Y(ttmp431),.A(g9941),.B(g9808));
OR2X1 OR_tmp432 (.Y(g9955),.A(g9947),.B(ttmp431));
OR2X1 OR_tmp433 (.Y(ttmp433),.A(g421),.B(I5576));
OR2X1 OR_tmp434 (.Y(ttmp434),.A(g448),.B(ttmp433));
OR2X1 OR_tmp435 (.Y(g2501),.A(g452),.B(ttmp434));
OR2X1 OR2_541 (.Y(g7231),.A(g6673),.B(g6087));
OR2X1 OR2_542 (.Y(g6078),.A(g4503),.B(g5256));
OR2X1 OR2_543 (.Y(g6478),.A(g5706),.B(g4967));
OR2X1 OR2_544 (.Y(g6907),.A(g6792),.B(g5675));
OR2X1 OR2_545 (.Y(g6035),.A(g5518),.B(g3974));
OR2X1 OR2_546 (.Y(g8937),.A(g8786),.B(g8698));
OR2X1 OR2_547 (.Y(g7742),.A(g7217),.B(g6743));
OR2X1 OR2_548 (.Y(g10722),.A(g10308),.B(g10671));
OR2X1 OR2_549 (.Y(g9918),.A(g9858),.B(g9698));
OR2X1 OR2_550 (.Y(g5403),.A(g4486),.B(g3695));
OR2X1 OR2_551 (.Y(g7926),.A(g7435),.B(g6892));
OR2X1 OR2_552 (.Y(g6915),.A(g6347),.B(g5686));
OR2X1 OR2_553 (.Y(g5841),.A(g4914),.B(g4230));
OR2X1 OR_tmp436 (.Y(ttmp436),.A(g9857),.B(g9877));
OR2X1 OR_tmp437 (.Y(ttmp437),.A(g9841),.B(ttmp436));
OR2X1 OR_tmp438 (.Y(I15220),.A(g9966),.B(ttmp437));
OR2X1 OR2_554 (.Y(g10529),.A(I16160),.B(I16161));
OR2X1 OR2_555 (.Y(g11246),.A(g11094),.B(g10948));
OR2X1 OR2_556 (.Y(g6002),.A(g5489),.B(g3939));
OR2X1 OR2_557 (.Y(g7712),.A(g7125),.B(g3540));
OR2X1 OR2_558 (.Y(g8810),.A(g7933),.B(g8720));
OR2X1 OR2_559 (.Y(g9921),.A(g9862),.B(g9703));
OR2X1 OR2_560 (.Y(g8432),.A(g8389),.B(g8072));
OR2X1 OR_tmp439 (.Y(ttmp439),.A(g9861),.B(g9874));
OR2X1 OR_tmp440 (.Y(ttmp440),.A(g9843),.B(ttmp439));
OR2X1 OR_tmp441 (.Y(I15172),.A(g9959),.B(ttmp440));
OR2X1 OR_tmp442 (.Y(ttmp442),.A(g9604),.B(g9582));
OR2X1 OR_tmp443 (.Y(I14822),.A(g9597),.B(ttmp442));
OR2X1 OR2_561 (.Y(g6928),.A(g6359),.B(g5703));
OR2X1 OR2_562 (.Y(g8157),.A(g7965),.B(g7623));
OR2X1 OR2_563 (.Y(g6930),.A(g6364),.B(g4269));
OR2X1 OR2_564 (.Y(g7660),.A(g7059),.B(g6583));
OR2X1 OR2_565 (.Y(g6899),.A(g6463),.B(g5471));
OR2X1 OR2_566 (.Y(g9392),.A(g9328),.B(g9324));
OR2X1 OR2_567 (.Y(g11318),.A(g11228),.B(g11104));
OR2X1 OR_tmp444 (.Y(ttmp444),.A(g10608),.B(g10604));
OR2X1 OR_tmp445 (.Y(I16427),.A(g10683),.B(ttmp444));
OR2X1 OR2_568 (.Y(g11227),.A(g11151),.B(g11010));
OR2X1 OR2_569 (.Y(g11058),.A(g10933),.B(g5280));
OR2X1 OR_tmp446 (.Y(ttmp446),.A(g1137),.B(g1133));
OR2X1 OR_tmp447 (.Y(ttmp447),.A(g1145),.B(ttmp446));
OR2X1 OR_tmp448 (.Y(I5351),.A(g1141),.B(ttmp447));
OR2X1 OR_tmp449 (.Y(ttmp449),.A(g9389),.B(g9646));
OR2X1 OR_tmp450 (.Y(g9708),.A(g9653),.B(ttmp449));
OR2X1 OR2_570 (.Y(g6071),.A(g5228),.B(g4505));
OR2X1 OR2_571 (.Y(g9911),.A(g9846),.B(g9689));
OR2X1 OR2_572 (.Y(g7102),.A(g6550),.B(g5915));
OR2X1 OR2_573 (.Y(g7302),.A(g7141),.B(g6328));
OR2X1 OR2_574 (.Y(g6038),.A(g5528),.B(g3979));
OR2X1 OR2_575 (.Y(g4239),.A(g4000),.B(g4008));
OR2X1 OR2_576 (.Y(g8646),.A(g8224),.B(g8547));
OR2X1 OR2_577 (.Y(g9974),.A(I15176),.B(I15177));
OR2X1 OR2_578 (.Y(g5823),.A(g5631),.B(g4882));
OR2X1 OR2_579 (.Y(g6918),.A(g6358),.B(g4252));
OR2X1 OR2_580 (.Y(g7265),.A(g6756),.B(g6204));
OR2X1 OR_tmp451 (.Y(ttmp451),.A(g2106),.B(g2104));
OR2X1 OR_tmp452 (.Y(ttmp452),.A(g2111),.B(ttmp451));
OR2X1 OR_tmp453 (.Y(I5804),.A(g2109),.B(ttmp452));
OR2X1 OR2_581 (.Y(g5851),.A(g4941),.B(g4253));
OR2X1 OR2_582 (.Y(g11481),.A(g6624),.B(g11458));
OR2X1 OR2_583 (.Y(g10336),.A(g10230),.B(g9572));
OR2X1 OR2_584 (.Y(g7296),.A(g7131),.B(g6322));
OR2X1 OR2_585 (.Y(g4300),.A(g3546),.B(g2391));
OR2X1 OR2_586 (.Y(g8647),.A(g8130),.B(g8470));
NAND2X1 NAND2_0 (.Y(g8546),.A(g3983),.B(g8390));
NAND2X1 NAND2_1 (.Y(g2516),.A(I5612),.B(I5613));
NAND2X1 NAND2_2 (.Y(g2987),.A(g2481),.B(g883));
NAND2X1 NAND2_3 (.Y(I5593),.A(g1703),.B(I5591));
NAND2X1 NAND2_4 (.Y(g8970),.A(g5548),.B(g8839));
NAND2X1 NAND2_5 (.Y(I10519),.A(g6231),.B(g822));
NAND2X1 NAND2_6 (.Y(I11279),.A(g305),.B(I11278));
AND2X1 AND_tmp454 (.Y(ttmp454),.A(g7562),.B(g7550));
AND2X1 AND_tmp455 (.Y(ttmp455),.A(g7011),.B(ttmp454));
NAND2X1 NAND_tmp456 (.Y(g7990),.A(g6995),.B(ttmp455));
NAND2X1 NAND2_7 (.Y(I11278),.A(g305),.B(g6485));
NAND2X1 NAND2_8 (.Y(g3978),.A(g3207),.B(g1822));
NAND2X1 NAND2_9 (.Y(I5264),.A(g456),.B(I5263));
NAND2X1 NAND2_10 (.Y(I8640),.A(g4278),.B(g516));
NAND2X1 NAND2_11 (.Y(I6761),.A(g2943),.B(I6760));
NAND2X1 NAND2_12 (.Y(I17400),.A(g11418),.B(g11416));
NAND2X1 NAND2_13 (.Y(I5450),.A(g1235),.B(I5449));
NAND2X1 NAND2_14 (.Y(I16060),.A(g10372),.B(I16058));
NAND2X1 NAND2_15 (.Y(I6746),.A(g2938),.B(g1453));
NAND2X1 NAND2_16 (.Y(I11975),.A(g1462),.B(I11973));
NAND2X1 NAND2_17 (.Y(I12136),.A(g7110),.B(g131));
NAND2X1 NAND2_18 (.Y(I11937),.A(g1458),.B(I11935));
NAND2X1 NAND2_19 (.Y(g2959),.A(I6167),.B(I6168));
NAND2X1 NAND2_20 (.Y(I5878),.A(g2120),.B(g2115));
NAND2X1 NAND2_21 (.Y(g2517),.A(I5619),.B(I5620));
NAND2X1 NAND2_22 (.Y(g5552),.A(g4777),.B(g4401));
NAND2X1 NAND2_23 (.Y(I6468),.A(g23),.B(I6467));
NAND2X1 NAND2_24 (.Y(I8796),.A(g4672),.B(I8795));
NAND2X1 NAND2_25 (.Y(g10392),.A(I15891),.B(I15892));
NAND2X1 NAND2_26 (.Y(I5611),.A(g1280),.B(g1284));
NAND2X1 NAND2_27 (.Y(g8738),.A(g8688),.B(g4921));
NAND2X1 NAND2_28 (.Y(I6716),.A(g201),.B(I6714));
NAND2X1 NAND2_29 (.Y(g2310),.A(g591),.B(g605));
NAND2X1 NAND2_30 (.Y(I7685),.A(g3460),.B(I7683));
NAND2X1 NAND2_31 (.Y(g3056),.A(g2374),.B(g599));
NAND2X1 NAND2_32 (.Y(I12108),.A(g135),.B(I12106));
AND2X1 AND_tmp457 (.Y(ttmp457),.A(g3062),.B(g2325));
NAND2X1 NAND_tmp458 (.Y(g3529),.A(g2310),.B(ttmp457));
NAND2X1 NAND2_33 (.Y(I6747),.A(g2938),.B(I6746));
NAND2X1 NAND2_34 (.Y(g2236),.A(I5230),.B(I5231));
NAND2X1 NAND2_35 (.Y(g7584),.A(I12075),.B(I12076));
NAND2X1 NAND2_36 (.Y(I15870),.A(g10358),.B(g2713));
NAND2X1 NAND2_37 (.Y(I16067),.A(g2765),.B(I16065));
NAND2X1 NAND2_38 (.Y(I7562),.A(g3533),.B(g654));
NAND2X1 NAND2_39 (.Y(I13531),.A(g8253),.B(I13529));
NAND2X1 NAND2_40 (.Y(I8797),.A(g1145),.B(I8795));
NAND2X1 NAND2_41 (.Y(I17584),.A(g11354),.B(g11515));
NAND2X1 NAND2_42 (.Y(I11936),.A(g7004),.B(I11935));
NAND2X1 NAND2_43 (.Y(I15257),.A(g9984),.B(I15256));
NAND2X1 NAND2_44 (.Y(g8402),.A(I13505),.B(I13506));
AND2X1 AND_tmp459 (.Y(ttmp459),.A(g8501),.B(g8739));
NAND2X1 NAND_tmp460 (.Y(g8824),.A(g8502),.B(ttmp459));
NAND2X1 NAND2_45 (.Y(I6186),.A(g2511),.B(g466));
NAND2X1 NAND2_46 (.Y(g11496),.A(I17504),.B(I17505));
NAND2X1 NAND2_47 (.Y(I16001),.A(g2683),.B(I15999));
NAND2X1 NAND2_48 (.Y(I6125),.A(g2215),.B(I6124));
NAND2X1 NAND2_49 (.Y(I11909),.A(g1474),.B(I11907));
NAND2X1 NAND2_50 (.Y(I12040),.A(g1466),.B(I12038));
NAND2X1 NAND2_51 (.Y(I13909),.A(g1432),.B(I13907));
NAND2X1 NAND2_52 (.Y(g3625),.A(I6771),.B(I6772));
NAND2X1 NAND2_53 (.Y(I11908),.A(g6967),.B(I11907));
NAND2X1 NAND2_54 (.Y(g10470),.A(I16008),.B(I16009));
NAND2X1 NAND2_55 (.Y(I13908),.A(g8526),.B(I13907));
NAND2X1 NAND2_56 (.Y(g3813),.A(I7034),.B(I7035));
NAND2X1 NAND2_57 (.Y(I8650),.A(g4824),.B(g778));
NAND2X1 NAND2_58 (.Y(g6207),.A(I9947),.B(I9948));
NAND2X1 NAND2_59 (.Y(I16066),.A(g10428),.B(I16065));
NAND2X1 NAND2_60 (.Y(g2948),.A(I6144),.B(I6145));
NAND2X1 NAND2_61 (.Y(I11242),.A(g6760),.B(I11241));
NAND2X1 NAND2_62 (.Y(g10467),.A(I15993),.B(I15994));
NAND2X1 NAND2_63 (.Y(I6187),.A(g2511),.B(I6186));
NAND2X1 NAND2_64 (.Y(g6488),.A(g6027),.B(g6019));
NAND2X1 NAND2_65 (.Y(I5500),.A(g1255),.B(g1007));
NAND2X1 NAND2_66 (.Y(I11974),.A(g7001),.B(I11973));
NAND2X1 NAND2_67 (.Y(I12062),.A(g1478),.B(I12060));
NAND2X1 NAND2_68 (.Y(g5300),.A(I8771),.B(I8772));
NAND2X1 NAND2_69 (.Y(I5184),.A(g1415),.B(g1515));
NAND2X1 NAND2_70 (.Y(I13293),.A(g1882),.B(g8161));
NAND2X1 NAND2_71 (.Y(I6200),.A(g2525),.B(I6199));
NAND2X1 NAND2_72 (.Y(I13265),.A(g1909),.B(g8154));
NAND2X1 NAND2_73 (.Y(I5024),.A(g995),.B(I5023));
NAND2X1 NAND2_74 (.Y(I7863),.A(g4099),.B(g774));
NAND2X1 NAND2_75 (.Y(g8705),.A(I13991),.B(I13992));
NAND2X1 NAND2_76 (.Y(g8471),.A(I13660),.B(I13661));
NAND2X1 NAND2_77 (.Y(I15256),.A(g9984),.B(g9980));
NAND2X1 NAND2_78 (.Y(I6145),.A(g646),.B(I6143));
NAND2X1 NAND2_79 (.Y(I13992),.A(g8688),.B(I13990));
NAND2X1 NAND2_80 (.Y(I11510),.A(g1806),.B(I11508));
NAND2X1 NAND2_81 (.Y(g10853),.A(g10731),.B(g5034));
NAND2X1 NAND2_82 (.Y(I5231),.A(g148),.B(I5229));
NAND2X1 NAND2_83 (.Y(I12047),.A(g1486),.B(I12045));
NAND2X1 NAND2_84 (.Y(I10771),.A(g1801),.B(I10769));
NAND2X1 NAND2_85 (.Y(g10477),.A(I16045),.B(I16046));
NAND2X1 NAND2_86 (.Y(g7582),.A(I12061),.B(I12062));
NAND2X1 NAND2_87 (.Y(I5104),.A(g431),.B(g435));
NAND2X1 NAND2_88 (.Y(g8409),.A(I13530),.B(I13531));
NAND2X1 NAND2_89 (.Y(I6447),.A(g2264),.B(g1776));
NAND2X1 NAND2_90 (.Y(I4956),.A(g327),.B(I4954));
NAND2X1 NAND2_91 (.Y(I5613),.A(g1284),.B(I5611));
NAND2X1 NAND2_92 (.Y(I8481),.A(g3530),.B(I8479));
NAND2X1 NAND2_93 (.Y(g5278),.A(I8739),.B(I8740));
NAND2X1 NAND2_94 (.Y(I6880),.A(g3301),.B(I6879));
NAND2X1 NAND2_95 (.Y(I15431),.A(g10047),.B(I15430));
NAND2X1 NAND2_96 (.Y(g5548),.A(g1840),.B(g4401));
AND2X1 AND_tmp461 (.Y(ttmp461),.A(g6984),.B(g6974));
AND2X1 AND_tmp462 (.Y(ttmp462),.A(g7011),.B(ttmp461));
NAND2X1 NAND_tmp463 (.Y(g7671),.A(g6995),.B(ttmp462));
NAND2X1 NAND2_97 (.Y(I12020),.A(g7119),.B(I12019));
NAND2X1 NAND2_98 (.Y(g10665),.A(I16331),.B(I16332));
NAND2X1 NAND2_99 (.Y(I16469),.A(g10518),.B(I16467));
NAND2X1 NAND2_100 (.Y(I5014),.A(g1007),.B(I5013));
NAND2X1 NAND2_101 (.Y(I13523),.A(g8249),.B(I13521));
NAND2X1 NAND2_102 (.Y(I16039),.A(g2707),.B(I16037));
NAND2X1 NAND2_103 (.Y(I16468),.A(g10716),.B(I16467));
NAND2X1 NAND2_104 (.Y(I12046),.A(g6951),.B(I12045));
NAND2X1 NAND2_105 (.Y(g4476),.A(g3807),.B(g3071));
NAND2X1 NAND2_106 (.Y(g10476),.A(I16038),.B(I16039));
NAND2X1 NAND2_107 (.Y(I16038),.A(g10427),.B(I16037));
NAND2X1 NAND2_108 (.Y(I8676),.A(g4374),.B(g1027));
NAND2X1 NAND2_109 (.Y(I12113),.A(g7093),.B(g162));
NAND2X1 NAND2_110 (.Y(I8761),.A(g4616),.B(g1129));
NAND2X1 NAND2_111 (.Y(g3204),.A(g2571),.B(g2061));
NAND2X1 NAND2_112 (.Y(I15993),.A(g10422),.B(I15992));
NAND2X1 NAND2_113 (.Y(I5036),.A(g1019),.B(I5034));
NAND2X1 NAND2_114 (.Y(I14263),.A(g8843),.B(g1814));
NAND2X1 NAND2_115 (.Y(g8298),.A(I13249),.B(I13250));
NAND2X1 NAND2_116 (.Y(I5135),.A(g521),.B(g525));
NAND2X1 NAND2_117 (.Y(g2405),.A(I5485),.B(I5486));
NAND2X1 NAND2_118 (.Y(I7034),.A(g3089),.B(I7033));
NAND2X1 NAND2_119 (.Y(I15443),.A(g10122),.B(I15441));
NAND2X1 NAND2_120 (.Y(I6166),.A(g2236),.B(g153));
NAND2X1 NAND2_121 (.Y(I8624),.A(g4267),.B(g511));
NAND2X1 NAND2_122 (.Y(I16015),.A(g10425),.B(g2695));
NAND2X1 NAND2_123 (.Y(I8677),.A(g4374),.B(I8676));
NAND2X1 NAND2_124 (.Y(I8576),.A(g4234),.B(I8575));
NAND2X1 NAND2_125 (.Y(I14613),.A(g9204),.B(I14612));
NAND2X1 NAND2_126 (.Y(I8716),.A(g4601),.B(I8715));
NAND2X1 NAND2_127 (.Y(g3530),.A(I6715),.B(I6716));
NAND2X1 NAND2_128 (.Y(g8405),.A(I13514),.B(I13515));
AND2X1 AND_tmp464 (.Y(ttmp464),.A(g2439),.B(g3200));
AND2X1 AND_tmp465 (.Y(ttmp465),.A(g3215),.B(ttmp464));
NAND2X1 NAND_tmp466 (.Y(g4104),.A(g3247),.B(ttmp465));
NAND2X1 NAND2_129 (.Y(I12003),.A(g7082),.B(I12002));
NAND2X1 NAND2_130 (.Y(g2177),.A(I5127),.B(I5128));
NAND2X1 NAND2_131 (.Y(g3010),.A(g2382),.B(g2399));
NAND2X1 NAND2_132 (.Y(g5179),.A(I8576),.B(I8577));
NAND2X1 NAND2_133 (.Y(I17395),.A(g11414),.B(I17393));
NAND2X1 NAND2_134 (.Y(g7067),.A(I11279),.B(I11280));
AND2X1 AND_tmp467 (.Y(ttmp467),.A(g6984),.B(g7550));
AND2X1 AND_tmp468 (.Y(ttmp468),.A(g7011),.B(ttmp467));
NAND2X1 NAND_tmp469 (.Y(g7994),.A(g7574),.B(ttmp468));
NAND2X1 NAND2_135 (.Y(I6167),.A(g2236),.B(I6166));
NAND2X1 NAND2_136 (.Y(I5265),.A(g461),.B(I5263));
NAND2X1 NAND2_137 (.Y(I6989),.A(g2760),.B(I6988));
NAND2X1 NAND2_138 (.Y(I13274),.A(g8158),.B(I13272));
NAND2X1 NAND2_139 (.Y(I10507),.A(g6221),.B(g786));
NAND2X1 NAND2_140 (.Y(I13530),.A(g704),.B(I13529));
NAND2X1 NAND2_141 (.Y(I5164),.A(g1508),.B(g1499));
NAND2X1 NAND2_142 (.Y(g9107),.A(I14443),.B(I14444));
NAND2X1 NAND2_143 (.Y(I9559),.A(g782),.B(I9557));
NAND2X1 NAND2_144 (.Y(I8577),.A(g496),.B(I8575));
NAND2X1 NAND2_145 (.Y(g2510),.A(I5592),.B(I5593));
NAND2X1 NAND2_146 (.Y(g8177),.A(I13077),.B(I13078));
NAND2X1 NAND2_147 (.Y(I8717),.A(g4052),.B(I8715));
NAND2X1 NAND2_148 (.Y(I5296),.A(g794),.B(I5295));
NAND2X1 NAND2_149 (.Y(g5209),.A(I8625),.B(I8626));
AND2X1 AND_tmp470 (.Y(ttmp470),.A(g7380),.B(g7273));
AND2X1 AND_tmp471 (.Y(ttmp471),.A(g7395),.B(ttmp470));
NAND2X1 NAND_tmp472 (.Y(g7950),.A(g7390),.B(ttmp471));
NAND2X1 NAND2_150 (.Y(g2088),.A(I4911),.B(I4912));
NAND2X1 NAND2_151 (.Y(I16000),.A(g10423),.B(I15999));
NAND2X1 NAND2_152 (.Y(I5371),.A(g971),.B(g976));
NAND2X1 NAND2_153 (.Y(g2215),.A(I5185),.B(I5186));
NAND2X1 NAND2_154 (.Y(g7101),.A(g6617),.B(g2364));
NAND2X1 NAND2_155 (.Y(I5675),.A(g1218),.B(g1223));
NAND2X1 NAND2_156 (.Y(I8544),.A(g4218),.B(I8543));
NAND2X1 NAND2_157 (.Y(g6577),.A(I10520),.B(I10521));
NAND2X1 NAND2_158 (.Y(I5297),.A(g798),.B(I5295));
NAND2X1 NAND2_159 (.Y(I13537),.A(g658),.B(g8157));
NAND2X1 NAND2_160 (.Y(I13283),.A(g1927),.B(g8159));
NAND2X1 NAND2_161 (.Y(g4749),.A(g3710),.B(g2061));
NAND2X1 NAND2_162 (.Y(I11982),.A(g1482),.B(I11980));
NAND2X1 NAND2_163 (.Y(I8514),.A(g4873),.B(I8513));
NAND2X1 NAND2_164 (.Y(I13091),.A(g1840),.B(I13089));
NAND2X1 NAND2_165 (.Y(g2943),.A(I6125),.B(I6126));
NAND2X1 NAND2_166 (.Y(I15908),.A(g10302),.B(I15906));
NAND2X1 NAND2_167 (.Y(I6879),.A(g3301),.B(g1351));
NAND2X1 NAND2_168 (.Y(I8763),.A(g1129),.B(I8761));
NAND2X1 NAND2_169 (.Y(I5449),.A(g1235),.B(g991));
AND2X1 AND_tmp473 (.Y(ttmp473),.A(g8738),.B(g8506));
NAND2X1 NAND_tmp474 (.Y(g8825),.A(g8502),.B(ttmp473));
NAND2X1 NAND2_170 (.Y(I16007),.A(g10424),.B(g2689));
NAND2X1 NAND2_171 (.Y(I5865),.A(g2107),.B(g2105));
NAND2X1 NAND2_172 (.Y(I5604),.A(g1149),.B(g1153));
NAND2X1 NAND2_173 (.Y(g2433),.A(I5517),.B(I5518));
NAND2X1 NAND2_174 (.Y(I6111),.A(g1494),.B(I6109));
NAND2X1 NAND2_175 (.Y(g2096),.A(I4929),.B(I4930));
NAND2X1 NAND2_176 (.Y(I13522),.A(g695),.B(I13521));
NAND2X1 NAND2_177 (.Y(I10770),.A(g5944),.B(I10769));
NAND2X1 NAND2_178 (.Y(g6027),.A(g4566),.B(g4921));
AND2X1 AND_tmp475 (.Y(ttmp475),.A(g6984),.B(g6974));
AND2X1 AND_tmp476 (.Y(ttmp476),.A(g7011),.B(ttmp475));
NAND2X1 NAND_tmp477 (.Y(g7992),.A(g7574),.B(ttmp476));
NAND2X1 NAND2_179 (.Y(I5539),.A(g1270),.B(I5538));
NAND2X1 NAND2_180 (.Y(I17394),.A(g11415),.B(I17393));
NAND2X1 NAND2_181 (.Y(I13553),.A(g668),.B(I13552));
NAND2X1 NAND2_182 (.Y(I8642),.A(g516),.B(I8640));
NAND2X1 NAND2_183 (.Y(g7573),.A(I12046),.B(I12047));
NAND2X1 NAND2_184 (.Y(g11416),.A(I17296),.B(I17297));
NAND2X1 NAND2_185 (.Y(g6003),.A(g5552),.B(g5548));
NAND2X1 NAND2_186 (.Y(g8934),.A(I14278),.B(I14279));
NAND2X1 NAND2_187 (.Y(I15992),.A(g10422),.B(g2677));
NAND2X1 NAND2_188 (.Y(I7683),.A(g1023),.B(g3460));
NAND2X1 NAND2_189 (.Y(I4910),.A(g386),.B(g318));
AND2X1 AND_tmp478 (.Y(ttmp478),.A(g2564),.B(g2571));
AND2X1 AND_tmp479 (.Y(ttmp479),.A(g2550),.B(ttmp478));
NAND2X1 NAND_tmp480 (.Y(g3209),.A(g2061),.B(ttmp479));
NAND2X1 NAND2_190 (.Y(I6794),.A(g143),.B(I6792));
NAND2X1 NAND2_191 (.Y(I10521),.A(g822),.B(I10519));
NAND2X1 NAND2_192 (.Y(I5486),.A(g1011),.B(I5484));
NAND2X1 NAND2_193 (.Y(I15442),.A(g10035),.B(I15441));
NAND2X1 NAND2_194 (.Y(g6858),.A(I10931),.B(I10932));
NAND2X1 NAND2_195 (.Y(I5185),.A(g1415),.B(I5184));
NAND2X1 NAND2_196 (.Y(g5304),.A(I8779),.B(I8780));
NAND2X1 NAND2_197 (.Y(g2354),.A(g1515),.B(g1520));
NAND2X1 NAND2_198 (.Y(I15615),.A(g10043),.B(g10153));
NAND2X1 NAND2_199 (.Y(I17281),.A(g11360),.B(g11357));
NAND2X1 NAND2_200 (.Y(I5470),.A(g999),.B(I5468));
NAND2X1 NAND2_201 (.Y(I11509),.A(g6580),.B(I11508));
NAND2X1 NAND2_202 (.Y(I5025),.A(g1275),.B(I5023));
NAND2X1 NAND2_203 (.Y(I11508),.A(g6580),.B(g1806));
NAND2X1 NAND2_204 (.Y(I15430),.A(g10047),.B(g10044));
NAND2X1 NAND2_205 (.Y(I14612),.A(g9204),.B(g611));
NAND2X1 NAND2_206 (.Y(g4675),.A(g4073),.B(g3247));
NAND2X1 NAND2_207 (.Y(I14272),.A(g1822),.B(I14270));
NAND2X1 NAND2_208 (.Y(g2979),.A(I6208),.B(I6209));
NAND2X1 NAND2_209 (.Y(I17290),.A(g11363),.B(I17288));
NAND2X1 NAND2_210 (.Y(g5269),.A(I8716),.B(I8717));
NAND2X1 NAND2_211 (.Y(g4297),.A(I7563),.B(I7564));
NAND2X1 NAND2_212 (.Y(I12002),.A(g7082),.B(g153));
NAND2X1 NAND2_213 (.Y(I5006),.A(g421),.B(I5005));
NAND2X1 NAND2_214 (.Y(I12128),.A(g170),.B(I12126));
NAND2X1 NAND2_215 (.Y(I5105),.A(g431),.B(I5104));
NAND2X1 NAND2_216 (.Y(I6323),.A(g2050),.B(I6322));
NAND2X1 NAND2_217 (.Y(g7588),.A(I12093),.B(I12094));
NAND2X1 NAND2_218 (.Y(I6666),.A(g2776),.B(I6664));
NAND2X1 NAND2_219 (.Y(g3623),.A(I6761),.B(I6762));
NAND2X1 NAND2_220 (.Y(I5373),.A(g976),.B(I5371));
NAND2X1 NAND2_221 (.Y(I8529),.A(g481),.B(I8527));
NAND2X1 NAND2_222 (.Y(I5283),.A(g758),.B(I5282));
NAND2X1 NAND2_223 (.Y(I7224),.A(g2981),.B(I7223));
NAND2X1 NAND2_224 (.Y(I5007),.A(g312),.B(I5005));
NAND2X1 NAND2_225 (.Y(I5459),.A(g1240),.B(g1003));
NAND2X1 NAND2_226 (.Y(I17297),.A(g11369),.B(I17295));
AND2X1 AND_tmp481 (.Y(ttmp481),.A(g6517),.B(g6509));
NAND2X1 NAND_tmp482 (.Y(g8746),.A(g8617),.B(ttmp481));
NAND2X1 NAND2_227 (.Y(I6143),.A(g1976),.B(g646));
NAND2X1 NAND2_228 (.Y(I5015),.A(g1011),.B(I5013));
NAND2X1 NAND2_229 (.Y(g8932),.A(I14264),.B(I14265));
NAND2X1 NAND2_230 (.Y(I16073),.A(g845),.B(I16072));
NAND2X1 NAND2_231 (.Y(I6988),.A(g2760),.B(g986));
NAND2X1 NAND2_232 (.Y(g3205),.A(g1814),.B(g2571));
NAND2X1 NAND2_233 (.Y(I8652),.A(g778),.B(I8650));
NAND2X1 NAND2_234 (.Y(I9558),.A(g5598),.B(I9557));
NAND2X1 NAND2_235 (.Y(I5203),.A(g369),.B(I5202));
NAND2X1 NAND2_236 (.Y(g7533),.A(I11936),.B(I11937));
NAND2X1 NAND2_237 (.Y(g3634),.A(I6806),.B(I6807));
NAND2X1 NAND2_238 (.Y(I6792),.A(g2959),.B(g143));
NAND2X1 NAND2_239 (.Y(g3304),.A(I6468),.B(I6469));
NAND2X1 NAND2_240 (.Y(I12145),.A(g158),.B(I12143));
NAND2X1 NAND2_241 (.Y(g7596),.A(I12127),.B(I12128));
NAND2X1 NAND2_242 (.Y(I13302),.A(g8162),.B(I13300));
NAND2X1 NAND2_243 (.Y(I5502),.A(g1007),.B(I5500));
NAND2X1 NAND2_244 (.Y(I9574),.A(g5608),.B(g818));
NAND2X1 NAND2_245 (.Y(g3273),.A(I6448),.B(I6449));
NAND2X1 NAND2_246 (.Y(I8670),.A(g4831),.B(I8669));
NAND2X1 NAND2_247 (.Y(I7035),.A(g1868),.B(I7033));
NAND2X1 NAND2_248 (.Y(I15453),.A(g10051),.B(I15451));
NAND2X1 NAND2_249 (.Y(I8625),.A(g4267),.B(I8624));
NAND2X1 NAND2_250 (.Y(I7876),.A(g4109),.B(I7875));
NAND2X1 NAND2_251 (.Y(I14203),.A(g8825),.B(I14202));
NAND2X1 NAND2_252 (.Y(I15607),.A(g10149),.B(g10144));
NAND2X1 NAND2_253 (.Y(g2274),.A(I5324),.B(I5325));
NAND2X1 NAND2_254 (.Y(I8740),.A(g1121),.B(I8738));
NAND2X1 NAND2_255 (.Y(I17296),.A(g11373),.B(I17295));
NAND2X1 NAND2_256 (.Y(g10507),.A(g10434),.B(g5859));
NAND2X1 NAND2_257 (.Y(g2325),.A(g611),.B(g617));
NAND2X1 NAND2_258 (.Y(I8606),.A(g506),.B(I8604));
NAND2X1 NAND2_259 (.Y(I12087),.A(g1470),.B(I12085));
NAND2X1 NAND2_260 (.Y(I13249),.A(g1891),.B(I13248));
NAND2X1 NAND2_261 (.Y(I13248),.A(g1891),.B(g8148));
NAND2X1 NAND2_262 (.Y(I13552),.A(g668),.B(g8262));
NAND2X1 NAND2_263 (.Y(g2106),.A(I4979),.B(I4980));
NAND2X1 NAND2_264 (.Y(I12069),.A(g139),.B(I12067));
NAND2X1 NAND2_265 (.Y(g9204),.A(g6019),.B(g8942));
NAND2X1 NAND2_266 (.Y(I12068),.A(g7116),.B(I12067));
NAND2X1 NAND2_267 (.Y(I17503),.A(g11475),.B(g7603));
NAND2X1 NAND2_268 (.Y(I7877),.A(g810),.B(I7875));
NAND2X1 NAND2_269 (.Y(I5165),.A(g1508),.B(I5164));
NAND2X1 NAND2_270 (.Y(g6740),.A(g6131),.B(g2550));
NAND2X1 NAND2_271 (.Y(I6289),.A(g981),.B(I6287));
NAND2X1 NAND2_272 (.Y(I6777),.A(g2892),.B(g650));
NAND2X1 NAND2_273 (.Y(g5171),.A(I8562),.B(I8563));
NAND2X1 NAND2_274 (.Y(I15891),.A(g853),.B(I15890));
NAND2X1 NAND2_275 (.Y(I13090),.A(g8006),.B(I13089));
NAND2X1 NAND2_276 (.Y(g11474),.A(I17460),.B(I17461));
AND2X1 AND_tmp483 (.Y(ttmp483),.A(g7380),.B(g7369));
AND2X1 AND_tmp484 (.Y(ttmp484),.A(g7395),.B(ttmp483));
NAND2X1 NAND_tmp485 (.Y(g7942),.A(g6847),.B(ttmp484));
NAND2X1 NAND2_277 (.Y(I5538),.A(g1270),.B(g1023));
NAND2X1 NAND2_278 (.Y(I7563),.A(g3533),.B(I7562));
NAND2X1 NAND2_279 (.Y(I13513),.A(g686),.B(g8248));
NAND2X1 NAND2_280 (.Y(g2107),.A(I4986),.B(I4987));
NAND2X1 NAND2_281 (.Y(g2223),.A(I5203),.B(I5204));
NAND2X1 NAND2_282 (.Y(I13505),.A(g677),.B(I13504));
NAND2X1 NAND2_283 (.Y(I6209),.A(g802),.B(I6207));
NAND2X1 NAND2_284 (.Y(I12086),.A(g6980),.B(I12085));
NAND2X1 NAND2_285 (.Y(I8545),.A(g486),.B(I8543));
NAND2X1 NAND2_286 (.Y(I8180),.A(g1786),.B(I8178));
NAND2X1 NAND2_287 (.Y(g2115),.A(I5014),.B(I5015));
NAND2X1 NAND2_288 (.Y(I8591),.A(g501),.B(I8589));
NAND2X1 NAND2_289 (.Y(I10931),.A(g6395),.B(I10930));
NAND2X1 NAND2_290 (.Y(I17402),.A(g11416),.B(I17400));
NAND2X1 NAND2_291 (.Y(g8307),.A(I13294),.B(I13295));
NAND2X1 NAND2_292 (.Y(I12144),.A(g7089),.B(I12143));
NAND2X1 NAND2_293 (.Y(I10520),.A(g6231),.B(I10519));
NAND2X1 NAND2_294 (.Y(I5263),.A(g456),.B(g461));
NAND2X1 NAND2_295 (.Y(g8757),.A(g8599),.B(g4401));
NAND2X1 NAND2_296 (.Y(I6714),.A(g2961),.B(g201));
NAND2X1 NAND2_297 (.Y(I14211),.A(g599),.B(I14209));
NAND2X1 NAND2_298 (.Y(I8515),.A(g3513),.B(I8513));
NAND2X1 NAND2_299 (.Y(g2272),.A(I5316),.B(I5317));
NAND2X1 NAND2_300 (.Y(I9946),.A(g5233),.B(g1796));
NAND2X1 NAND2_301 (.Y(I8750),.A(g4613),.B(g1125));
NAND2X1 NAND2_302 (.Y(I5605),.A(g1149),.B(I5604));
NAND2X1 NAND2_303 (.Y(g8880),.A(I14203),.B(I14204));
NAND2X1 NAND2_304 (.Y(I16051),.A(g837),.B(g10371));
NAND2X1 NAND2_305 (.Y(I16072),.A(g845),.B(g10373));
NAND2X1 NAND2_306 (.Y(g10440),.A(g10360),.B(g6037));
NAND2X1 NAND2_307 (.Y(g8612),.A(I13858),.B(I13859));
NAND2X1 NAND2_308 (.Y(I15872),.A(g2713),.B(I15870));
NAND2X1 NAND2_309 (.Y(I8528),.A(g4879),.B(I8527));
NAND2X1 NAND2_310 (.Y(g8629),.A(I13901),.B(I13902));
AND2X1 AND_tmp486 (.Y(ttmp486),.A(g1814),.B(g8390));
AND2X1 AND_tmp487 (.Y(ttmp487),.A(g2571),.B(ttmp486));
NAND2X1 NAND_tmp488 (.Y(g8542),.A(g1828),.B(ttmp487));
NAND2X1 NAND2_311 (.Y(I9947),.A(g5233),.B(I9946));
NAND2X1 NAND2_312 (.Y(I6838),.A(g806),.B(I6836));
NAND2X1 NAND2_313 (.Y(g7583),.A(I12068),.B(I12069));
NAND2X1 NAND2_314 (.Y(g4803),.A(g3664),.B(g2356));
NAND2X1 NAND2_315 (.Y(I17307),.A(g11377),.B(I17305));
NAND2X1 NAND2_316 (.Y(g4538),.A(g3475),.B(g2399));
NAND2X1 NAND2_317 (.Y(I15452),.A(g10058),.B(I15451));
NAND2X1 NAND2_318 (.Y(I13857),.A(g8538),.B(g1448));
NAND2X1 NAND2_319 (.Y(I14202),.A(g8825),.B(g591));
NAND2X1 NAND2_320 (.Y(I13765),.A(g731),.B(g8417));
NAND2X1 NAND2_321 (.Y(g2260),.A(I5296),.B(I5297));
AND2X1 AND_tmp489 (.Y(ttmp489),.A(g6984),.B(g7550));
AND2X1 AND_tmp490 (.Y(ttmp490),.A(g7011),.B(ttmp489));
NAND2X1 NAND_tmp491 (.Y(g7986),.A(g6995),.B(ttmp490));
NAND2X1 NAND2_322 (.Y(g5226),.A(I8670),.B(I8671));
NAND2X1 NAND2_323 (.Y(g8512),.A(g3723),.B(g8366));
NAND2X1 NAND2_324 (.Y(I16046),.A(g10370),.B(I16044));
NAND2X1 NAND2_325 (.Y(I13504),.A(g677),.B(g8247));
NAND2X1 NAND2_326 (.Y(g10447),.A(g10363),.B(g5360));
NAND2X1 NAND2_327 (.Y(g2167),.A(I5105),.B(I5106));
NAND2X1 NAND2_328 (.Y(I8804),.A(g4677),.B(I8803));
NAND2X1 NAND2_329 (.Y(g10472),.A(I16016),.B(I16017));
NAND2X1 NAND2_330 (.Y(I17487),.A(g11474),.B(I17485));
NAND2X1 NAND2_331 (.Y(I4995),.A(g416),.B(g309));
NAND2X1 NAND2_332 (.Y(I12093),.A(g6944),.B(I12092));
AND2X1 AND_tmp492 (.Y(ttmp492),.A(g7562),.B(g6974));
AND2X1 AND_tmp493 (.Y(ttmp493),.A(g7011),.B(ttmp492));
NAND2X1 NAND_tmp494 (.Y(g7987),.A(g6995),.B(ttmp493));
NAND2X1 NAND2_333 (.Y(g5227),.A(I8677),.B(I8678));
NAND2X1 NAND2_334 (.Y(I5126),.A(g1386),.B(g1389));
NAND2X1 NAND2_335 (.Y(g2321),.A(I5372),.B(I5373));
NAND2X1 NAND2_336 (.Y(g7547),.A(I11974),.B(I11975));
NAND2X1 NAND2_337 (.Y(I17306),.A(g11381),.B(I17305));
AND2X1 AND_tmp495 (.Y(ttmp495),.A(g6124),.B(g6122));
NAND2X1 NAND_tmp496 (.Y(g6548),.A(g6132),.B(ttmp495));
NAND2X1 NAND2_338 (.Y(I11995),.A(g7107),.B(g127));
NAND2X1 NAND2_339 (.Y(I7225),.A(g1781),.B(I7223));
NAND2X1 NAND2_340 (.Y(I11261),.A(g6775),.B(g826));
AND2X1 AND_tmp497 (.Y(ttmp497),.A(g8757),.B(g8545));
NAND2X1 NAND_tmp498 (.Y(g8843),.A(g8542),.B(ttmp497));
NAND2X1 NAND2_341 (.Y(g2938),.A(I6110),.B(I6111));
NAND2X1 NAND2_342 (.Y(I4942),.A(g396),.B(I4941));
NAND2X1 NAND2_343 (.Y(g10394),.A(I15899),.B(I15900));
NAND2X1 NAND2_344 (.Y(g8549),.A(g5527),.B(g8390));
NAND2X1 NAND2_345 (.Y(g3070),.A(g2016),.B(g1206));
NAND2X1 NAND2_346 (.Y(I4954),.A(g401),.B(g327));
NAND2X1 NAND2_347 (.Y(I5023),.A(g995),.B(g1275));
NAND2X1 NAND2_348 (.Y(g10446),.A(g10443),.B(g5350));
NAND2X1 NAND2_349 (.Y(I16081),.A(g10374),.B(I16079));
NAND2X1 NAND2_350 (.Y(I8641),.A(g4278),.B(I8640));
NAND2X1 NAND2_351 (.Y(I6178),.A(g197),.B(I6176));
NAND2X1 NAND2_352 (.Y(I12075),.A(g7098),.B(I12074));
NAND2X1 NAND2_353 (.Y(I5127),.A(g1386),.B(I5126));
NAND2X1 NAND2_354 (.Y(I5451),.A(g991),.B(I5449));
NAND2X1 NAND2_355 (.Y(g4168),.A(I7322),.B(I7323));
NAND2X1 NAND2_356 (.Y(I6288),.A(g2091),.B(I6287));
NAND2X1 NAND2_357 (.Y(I8179),.A(g3685),.B(I8178));
NAND2X1 NAND2_358 (.Y(I4912),.A(g318),.B(I4910));
NAND2X1 NAND2_359 (.Y(I6805),.A(g3268),.B(g471));
AND2X1 AND_tmp499 (.Y(ttmp499),.A(g3222),.B(g2493));
NAND2X1 NAND_tmp500 (.Y(g3766),.A(g2439),.B(ttmp499));
NAND2X1 NAND2_360 (.Y(g3087),.A(I6288),.B(I6289));
NAND2X1 NAND2_361 (.Y(I17486),.A(g11384),.B(I17485));
NAND2X1 NAND2_362 (.Y(I4929),.A(g391),.B(I4928));
NAND2X1 NAND2_363 (.Y(I15890),.A(g853),.B(g10286));
NAND2X1 NAND2_364 (.Y(I16331),.A(g10616),.B(I16330));
NAND2X1 NAND2_365 (.Y(I9575),.A(g5608),.B(I9574));
NAND2X1 NAND2_366 (.Y(I13887),.A(g8532),.B(I13886));
NAND2X1 NAND2_367 (.Y(g5308),.A(I8787),.B(I8788));
NAND2X1 NAND2_368 (.Y(I13529),.A(g704),.B(g8253));
NAND2X1 NAND2_369 (.Y(I6208),.A(g2534),.B(I6207));
NAND2X1 NAND2_370 (.Y(g5217),.A(I8641),.B(I8642));
NAND2X1 NAND2_371 (.Y(I5316),.A(g1032),.B(I5315));
NAND2X1 NAND2_372 (.Y(g2111),.A(I5006),.B(I5007));
NAND2X1 NAND2_373 (.Y(g10366),.A(g10285),.B(g5392));
NAND2X1 NAND2_374 (.Y(I5034),.A(g1015),.B(g1019));
NAND2X1 NAND2_375 (.Y(I13869),.A(g1403),.B(I13867));
NAND2X1 NAND2_376 (.Y(I13868),.A(g8523),.B(I13867));
NAND2X1 NAND2_377 (.Y(I15999),.A(g10423),.B(g2683));
NAND2X1 NAND2_378 (.Y(I13259),.A(g1900),.B(I13258));
AND2X1 AND_tmp501 (.Y(ttmp501),.A(g2211),.B(g2202));
AND2X1 AND_tmp502 (.Y(ttmp502),.A(g2229),.B(ttmp501));
NAND2X1 NAND_tmp503 (.Y(g3261),.A(g2222),.B(ttmp502));
NAND2X1 NAND2_379 (.Y(g10481),.A(I16073),.B(I16074));
NAND2X1 NAND2_380 (.Y(g2180),.A(I5136),.B(I5137));
AND2X1 AND_tmp504 (.Y(ttmp504),.A(g4604),.B(g3807));
NAND2X1 NAND_tmp505 (.Y(g4976),.A(g2310),.B(ttmp504));
NAND2X1 NAND2_381 (.Y(g8506),.A(g3475),.B(g8366));
NAND2X1 NAND2_382 (.Y(g2380),.A(I5460),.B(I5461));
NAND2X1 NAND2_383 (.Y(I13258),.A(g1900),.B(g8153));
NAND2X1 NAND2_384 (.Y(I5013),.A(g1007),.B(g1011));
NAND2X1 NAND2_385 (.Y(g5196),.A(I8605),.B(I8606));
NAND2X1 NAND2_386 (.Y(I10930),.A(g6395),.B(g5555));
NAND2X1 NAND2_387 (.Y(I6770),.A(g3257),.B(g382));
NAND2X1 NAND2_388 (.Y(g11449),.A(I17401),.B(I17402));
NAND2X1 NAND2_389 (.Y(g11448),.A(I17394),.B(I17395));
NAND2X1 NAND2_390 (.Y(I15717),.A(g10231),.B(I15716));
NAND2X1 NAND2_391 (.Y(I5317),.A(g1027),.B(I5315));
NAND2X1 NAND2_392 (.Y(I14210),.A(g8824),.B(I14209));
NAND2X1 NAND2_393 (.Y(I17569),.A(g1610),.B(I17567));
NAND2X1 NAND2_394 (.Y(I13878),.A(g1444),.B(I13876));
NAND2X1 NAND2_395 (.Y(g8545),.A(g3710),.B(g8390));
NAND2X1 NAND2_396 (.Y(g2515),.A(I5605),.B(I5606));
NAND2X1 NAND2_397 (.Y(I14443),.A(g8970),.B(I14442));
NAND2X1 NAND2_398 (.Y(g7557),.A(I11996),.B(I11997));
NAND2X1 NAND2_399 (.Y(g8180),.A(I13090),.B(I13091));
NAND2X1 NAND2_400 (.Y(I14279),.A(g1828),.B(I14277));
NAND2X1 NAND2_401 (.Y(I17568),.A(g11496),.B(I17567));
NAND2X1 NAND2_402 (.Y(I13886),.A(g8532),.B(g1440));
NAND2X1 NAND2_403 (.Y(I7322),.A(g3047),.B(I7321));
NAND2X1 NAND2_404 (.Y(I6990),.A(g986),.B(I6988));
NAND2X1 NAND2_405 (.Y(I14278),.A(g8847),.B(I14277));
NAND2X1 NAND2_406 (.Y(I7033),.A(g3089),.B(g1868));
NAND2X1 NAND2_407 (.Y(I9006),.A(g4492),.B(g1791));
NAND2X1 NAND2_408 (.Y(g8507),.A(g3738),.B(g8366));
NAND2X1 NAND2_409 (.Y(I5460),.A(g1240),.B(I5459));
NAND2X1 NAND2_410 (.Y(g4588),.A(g3440),.B(g2745));
NAND2X1 NAND2_411 (.Y(I4986),.A(g999),.B(I4985));
AND2X1 AND_tmp506 (.Y(ttmp506),.A(g2564),.B(g2571));
NAND2X1 NAND_tmp507 (.Y(g3247),.A(g1828),.B(ttmp506));
NAND2X1 NAND2_412 (.Y(I8651),.A(g4824),.B(I8650));
NAND2X1 NAND2_413 (.Y(I13545),.A(g713),.B(I13544));
NAND2X1 NAND2_414 (.Y(g8628),.A(I13894),.B(I13895));
NAND2X1 NAND2_415 (.Y(I6138),.A(g378),.B(I6136));
NAND2X1 NAND2_416 (.Y(I12074),.A(g7098),.B(g174));
NAND2X1 NAND2_417 (.Y(g8630),.A(I13908),.B(I13909));
NAND2X1 NAND2_418 (.Y(I13078),.A(g7963),.B(I13076));
NAND2X1 NAND2_419 (.Y(I6109),.A(g2205),.B(g1494));
NAND2X1 NAND2_420 (.Y(g8300),.A(I13259),.B(I13260));
NAND2X1 NAND2_421 (.Y(I5501),.A(g1255),.B(I5500));
NAND2X1 NAND2_422 (.Y(I17586),.A(g11515),.B(I17584));
NAND2X1 NAND2_423 (.Y(I12092),.A(g6944),.B(g1490));
NAND2X1 NAND2_424 (.Y(I13901),.A(g8520),.B(I13900));
NAND2X1 NAND2_425 (.Y(I8795),.A(g4672),.B(g1145));
NAND2X1 NAND2_426 (.Y(I6201),.A(g766),.B(I6199));
NAND2X1 NAND2_427 (.Y(I14217),.A(g8826),.B(I14216));
NAND2X1 NAND2_428 (.Y(I9007),.A(g4492),.B(I9006));
NAND2X1 NAND2_429 (.Y(I13561),.A(g8263),.B(I13559));
NAND2X1 NAND2_430 (.Y(I15716),.A(g10231),.B(g10229));
NAND2X1 NAND2_431 (.Y(I6449),.A(g1776),.B(I6447));
NAND2X1 NAND2_432 (.Y(I13295),.A(g8161),.B(I13293));
NAND2X1 NAND2_433 (.Y(I4987),.A(g1003),.B(I4985));
NAND2X1 NAND2_434 (.Y(I6715),.A(g2961),.B(I6714));
NAND2X1 NAND2_435 (.Y(I17493),.A(g11475),.B(I17492));
NAND2X1 NAND2_436 (.Y(I12215),.A(g7061),.B(I12214));
NAND2X1 NAND2_437 (.Y(g2372),.A(I5450),.B(I5451));
NAND2X1 NAND2_438 (.Y(g7062),.A(I11262),.B(I11263));
NAND2X1 NAND2_439 (.Y(g2988),.A(I6225),.B(I6226));
NAND2X1 NAND2_440 (.Y(I13309),.A(g617),.B(I13307));
NAND2X1 NAND2_441 (.Y(g8839),.A(g8750),.B(g4401));
NAND2X1 NAND2_442 (.Y(g2555),.A(I5676),.B(I5677));
NAND2X1 NAND2_443 (.Y(g3662),.A(I6826),.B(I6827));
NAND2X1 NAND2_444 (.Y(I13308),.A(g8190),.B(I13307));
NAND2X1 NAND2_445 (.Y(g2792),.A(I5879),.B(I5880));
NAND2X1 NAND2_446 (.Y(g4117),.A(g3041),.B(g3061));
NAND2X1 NAND2_447 (.Y(I8543),.A(g4218),.B(g486));
NAND2X1 NAND2_448 (.Y(g11549),.A(I17585),.B(I17586));
NAND2X1 NAND2_449 (.Y(I6881),.A(g1351),.B(I6879));
NAND2X1 NAND2_450 (.Y(I12138),.A(g131),.B(I12136));
NAND2X1 NAND2_451 (.Y(I8729),.A(g4605),.B(I8728));
NAND2X1 NAND2_452 (.Y(I14216),.A(g8826),.B(g605));
NAND2X1 NAND2_453 (.Y(g10384),.A(I15871),.B(I15872));
NAND2X1 NAND2_454 (.Y(I13260),.A(g8153),.B(I13258));
NAND2X1 NAND2_455 (.Y(g2776),.A(I5866),.B(I5867));
NAND2X1 NAND2_456 (.Y(I8513),.A(g4873),.B(g3513));
NAND2X1 NAND2_457 (.Y(I13559),.A(g722),.B(g8263));
NAND2X1 NAND2_458 (.Y(I8178),.A(g3685),.B(g1786));
NAND2X1 NAND2_459 (.Y(g3631),.A(I6793),.B(I6794));
NAND2X1 NAND2_460 (.Y(I6487),.A(g2306),.B(g1227));
NAND2X1 NAND2_461 (.Y(I16080),.A(g849),.B(I16079));
NAND2X1 NAND2_462 (.Y(I13893),.A(g8529),.B(g1436));
NAND2X1 NAND2_463 (.Y(I12115),.A(g162),.B(I12113));
NAND2X1 NAND2_464 (.Y(I6748),.A(g1453),.B(I6746));
NAND2X1 NAND2_465 (.Y(I13544),.A(g713),.B(g8259));
NAND2X1 NAND2_466 (.Y(I5484),.A(g1250),.B(g1011));
NAND2X1 NAND2_467 (.Y(I4928),.A(g391),.B(g321));
NAND2X1 NAND2_468 (.Y(I6226),.A(g1346),.B(I6224));
NAND2X1 NAND2_469 (.Y(I8805),.A(g1113),.B(I8803));
NAND2X1 NAND2_470 (.Y(I4930),.A(g321),.B(I4928));
NAND2X1 NAND2_471 (.Y(I15880),.A(g2719),.B(I15878));
NAND2X1 NAND2_472 (.Y(I14265),.A(g1814),.B(I14263));
NAND2X1 NAND2_473 (.Y(I16031),.A(g829),.B(I16030));
NAND2X1 NAND2_474 (.Y(g3585),.A(I6747),.B(I6748));
AND2X1 AND_tmp508 (.Y(ttmp508),.A(g2374),.B(g2382));
AND2X1 AND_tmp509 (.Y(ttmp509),.A(g2364),.B(ttmp508));
NAND2X1 NAND_tmp510 (.Y(g3041),.A(g2399),.B(ttmp509));
NAND2X1 NAND2_475 (.Y(g8933),.A(I14271),.B(I14272));
NAND2X1 NAND2_476 (.Y(I16330),.A(g10616),.B(g4997));
NAND2X1 NAND2_477 (.Y(I13267),.A(g8154),.B(I13265));
NAND2X1 NAND2_478 (.Y(I13294),.A(g1882),.B(I13293));
NAND2X1 NAND2_479 (.Y(g10231),.A(I15616),.B(I15617));
NAND2X1 NAND2_480 (.Y(I14442),.A(g8970),.B(g1834));
NAND2X1 NAND2_481 (.Y(I6793),.A(g2959),.B(I6792));
NAND2X1 NAND2_482 (.Y(I4966),.A(g330),.B(I4964));
NAND2X1 NAND2_483 (.Y(I8752),.A(g1125),.B(I8750));
NAND2X1 NAND2_484 (.Y(I15432),.A(g10044),.B(I15430));
NAND2X1 NAND2_485 (.Y(I12214),.A(g7061),.B(g2518));
NAND2X1 NAND2_486 (.Y(g10511),.A(g10438),.B(g6032));
NAND2X1 NAND2_487 (.Y(g3011),.A(g591),.B(g2382));
NAND2X1 NAND2_488 (.Y(g5103),.A(I8480),.B(I8481));
NAND2X1 NAND2_489 (.Y(I16087),.A(g861),.B(I16086));
NAND2X1 NAND2_490 (.Y(g3734),.A(g3039),.B(g599));
NAND2X1 NAND2_491 (.Y(I6664),.A(g2792),.B(g2776));
NAND2X1 NAND2_492 (.Y(g8882),.A(I14217),.B(I14218));
NAND2X1 NAND2_493 (.Y(I4955),.A(g401),.B(I4954));
NAND2X1 NAND2_494 (.Y(I8786),.A(g4639),.B(g1141));
AND2X1 AND_tmp511 (.Y(ttmp511),.A(g2550),.B(g2990));
NAND2X1 NAND_tmp512 (.Y(g3992),.A(g2571),.B(ttmp511));
NAND2X1 NAND2_495 (.Y(g10480),.A(I16066),.B(I16067));
NAND2X1 NAND2_496 (.Y(I11915),.A(g6935),.B(I11914));
NAND2X1 NAND2_497 (.Y(I8770),.A(g4619),.B(g1133));
NAND2X1 NAND2_498 (.Y(I5516),.A(g1260),.B(g1019));
NAND2X1 NAND2_499 (.Y(g8541),.A(g4001),.B(g8390));
NAND2X1 NAND2_500 (.Y(I6188),.A(g466),.B(I6186));
NAND2X1 NAND2_501 (.Y(g5147),.A(I8544),.B(I8545));
AND2X1 AND_tmp513 (.Y(ttmp513),.A(g6509),.B(g6971));
NAND2X1 NAND_tmp514 (.Y(g8744),.A(g8617),.B(ttmp513));
NAND2X1 NAND2_502 (.Y(I5892),.A(g750),.B(I5891));
NAND2X1 NAND2_503 (.Y(g8558),.A(I13766),.B(I13767));
NAND2X1 NAND2_504 (.Y(I15258),.A(g9980),.B(I15256));
NAND2X1 NAND2_505 (.Y(I13266),.A(g1909),.B(I13265));
NAND2X1 NAND2_506 (.Y(I8787),.A(g4639),.B(I8786));
NAND2X1 NAND2_507 (.Y(I6826),.A(g3281),.B(I6825));
NAND2X1 NAND2_508 (.Y(I17283),.A(g11357),.B(I17281));
AND2X1 AND_tmp515 (.Y(ttmp515),.A(g3247),.B(g3205));
NAND2X1 NAND_tmp516 (.Y(g5013),.A(g4749),.B(ttmp515));
NAND2X1 NAND2_509 (.Y(I17492),.A(g11475),.B(g3623));
NAND2X1 NAND2_510 (.Y(g8511),.A(g5277),.B(g8366));
NAND2X1 NAND2_511 (.Y(I16079),.A(g849),.B(g10374));
NAND2X1 NAND2_512 (.Y(I5035),.A(g1015),.B(I5034));
NAND2X1 NAND2_513 (.Y(I5517),.A(g1260),.B(I5516));
NAND2X1 NAND2_514 (.Y(I7223),.A(g2981),.B(g1781));
NAND2X1 NAND2_515 (.Y(I16086),.A(g861),.B(g10375));
NAND2X1 NAND2_516 (.Y(g5317),.A(I8796),.B(I8797));
NAND2X1 NAND2_517 (.Y(I15879),.A(g10359),.B(I15878));
NAND2X1 NAND2_518 (.Y(I15878),.A(g10359),.B(g2719));
NAND2X1 NAND2_519 (.Y(I12114),.A(g7093),.B(I12113));
NAND2X1 NAND2_520 (.Y(I12107),.A(g7113),.B(I12106));
NAND2X1 NAND2_521 (.Y(g2500),.A(g178),.B(g182));
NAND2X1 NAND2_522 (.Y(I15994),.A(g2677),.B(I15992));
AND2X1 AND_tmp517 (.Y(ttmp517),.A(g7279),.B(g7369));
AND2X1 AND_tmp518 (.Y(ttmp518),.A(g7395),.B(ttmp517));
NAND2X1 NAND_tmp519 (.Y(g7934),.A(g6847),.B(ttmp518));
NAND2X1 NAND2_523 (.Y(g10469),.A(g10430),.B(g5999));
NAND2X1 NAND2_524 (.Y(I14264),.A(g8843),.B(I14263));
NAND2X1 NAND2_525 (.Y(I6448),.A(g2264),.B(I6447));
NAND2X1 NAND2_526 (.Y(I13285),.A(g8159),.B(I13283));
NAND2X1 NAND2_527 (.Y(g10468),.A(I16000),.B(I16001));
NAND2X1 NAND2_528 (.Y(I6827),.A(g770),.B(I6825));
NAND2X1 NAND2_529 (.Y(g8623),.A(I13877),.B(I13878));
NAND2X1 NAND2_530 (.Y(I13900),.A(g8520),.B(g1428));
NAND2X1 NAND2_531 (.Y(g2795),.A(I5892),.B(I5893));
NAND2X1 NAND2_532 (.Y(I8575),.A(g4234),.B(g496));
NAND2X1 NAND2_533 (.Y(I14209),.A(g8824),.B(g599));
NAND2X1 NAND2_534 (.Y(I13560),.A(g722),.B(I13559));
NAND2X1 NAND2_535 (.Y(I8715),.A(g4601),.B(g4052));
NAND2X1 NAND2_536 (.Y(I8604),.A(g4259),.B(g506));
NAND2X1 NAND2_537 (.Y(I16017),.A(g2695),.B(I16015));
NAND2X1 NAND2_538 (.Y(I4941),.A(g396),.B(g324));
NAND2X1 NAND2_539 (.Y(g2205),.A(I5165),.B(I5166));
AND2X1 AND_tmp520 (.Y(ttmp520),.A(g2364),.B(g2800));
NAND2X1 NAND_tmp521 (.Y(g3753),.A(g2382),.B(ttmp520));
NAND2X1 NAND2_540 (.Y(I6467),.A(g23),.B(g2479));
NAND2X1 NAND2_541 (.Y(I14614),.A(g611),.B(I14612));
NAND2X1 NAND2_542 (.Y(g2104),.A(I4965),.B(I4966));
NAND2X1 NAND2_543 (.Y(g2099),.A(I4942),.B(I4943));
NAND2X1 NAND2_544 (.Y(I16023),.A(g10426),.B(g2701));
NAND2X1 NAND2_545 (.Y(g10479),.A(I16059),.B(I16060));
AND2X1 AND_tmp522 (.Y(ttmp522),.A(g4921),.B(g8688));
NAND2X1 NAND_tmp523 (.Y(g8737),.A(g2317),.B(ttmp522));
NAND2X1 NAND2_546 (.Y(g5942),.A(I9575),.B(I9576));
NAND2X1 NAND2_547 (.Y(g10478),.A(I16052),.B(I16053));
NAND2X1 NAND2_548 (.Y(I12004),.A(g153),.B(I12002));
NAND2X1 NAND2_549 (.Y(I4911),.A(g386),.B(I4910));
NAND2X1 NAND2_550 (.Y(I11914),.A(g6935),.B(g1494));
NAND2X1 NAND2_551 (.Y(g7960),.A(g7409),.B(g5573));
NAND2X1 NAND2_552 (.Y(I5295),.A(g794),.B(g798));
NAND2X1 NAND2_553 (.Y(I12106),.A(g7113),.B(g135));
NAND2X1 NAND2_554 (.Y(I8728),.A(g4605),.B(g1117));
NAND2X1 NAND2_555 (.Y(g3681),.A(I6837),.B(I6838));
NAND2X1 NAND2_556 (.Y(I11907),.A(g6967),.B(g1474));
NAND2X1 NAND2_557 (.Y(I13907),.A(g8526),.B(g1432));
NAND2X1 NAND2_558 (.Y(I8730),.A(g1117),.B(I8728));
NAND2X1 NAND2_559 (.Y(g8551),.A(g3967),.B(g8390));
NAND2X1 NAND2_560 (.Y(I4980),.A(g333),.B(I4978));
NAND2X1 NAND2_561 (.Y(g2961),.A(I6177),.B(I6178));
NAND2X1 NAND2_562 (.Y(g6019),.A(g617),.B(g4921));
NAND2X1 NAND2_563 (.Y(I16016),.A(g10425),.B(I16015));
NAND2X1 NAND2_564 (.Y(I11935),.A(g7004),.B(g1458));
NAND2X1 NAND2_565 (.Y(I8678),.A(g1027),.B(I8676));
NAND2X1 NAND2_566 (.Y(I17051),.A(g10923),.B(g11249));
NAND2X1 NAND2_567 (.Y(g4482),.A(I7864),.B(I7865));
NAND2X1 NAND2_568 (.Y(g7592),.A(I12107),.B(I12108));
NAND2X1 NAND2_569 (.Y(g3460),.A(I6665),.B(I6666));
AND2X1 AND_tmp524 (.Y(ttmp524),.A(g7279),.B(g7273));
AND2X1 AND_tmp525 (.Y(ttmp525),.A(g7395),.B(ttmp524));
NAND2X1 NAND_tmp526 (.Y(g7932),.A(g6847),.B(ttmp525));
NAND2X1 NAND2_570 (.Y(g7624),.A(I12215),.B(I12216));
AND2X1 AND_tmp527 (.Y(ttmp527),.A(g7380),.B(g7369));
AND2X1 AND_tmp528 (.Y(ttmp528),.A(g7395),.B(ttmp527));
NAND2X1 NAND_tmp529 (.Y(g7953),.A(g7390),.B(ttmp528));
NAND2X1 NAND2_571 (.Y(g8414),.A(I13553),.B(I13554));
NAND2X1 NAND2_572 (.Y(I6168),.A(g153),.B(I6166));
NAND2X1 NAND2_573 (.Y(I5229),.A(g182),.B(g148));
NAND2X1 NAND2_574 (.Y(I6772),.A(g382),.B(I6770));
NAND2X1 NAND2_575 (.Y(I16030),.A(g829),.B(g10368));
NAND2X1 NAND2_576 (.Y(I13284),.A(g1927),.B(I13283));
NAND2X1 NAND2_577 (.Y(I16065),.A(g10428),.B(g2765));
NAND2X1 NAND2_578 (.Y(g2947),.A(I6137),.B(I6138));
NAND2X1 NAND2_579 (.Y(I7321),.A(g3047),.B(g1231));
NAND2X1 NAND2_580 (.Y(g2437),.A(I5529),.B(I5530));
NAND2X1 NAND2_581 (.Y(g2102),.A(I4955),.B(I4956));
NAND2X1 NAND2_582 (.Y(I17282),.A(g11360),.B(I17281));
NAND2X1 NAND2_583 (.Y(I5620),.A(g1771),.B(I5618));
NAND2X1 NAND2_584 (.Y(I8664),.A(g476),.B(I8662));
NAND2X1 NAND2_585 (.Y(g7524),.A(I11915),.B(I11916));
NAND2X1 NAND2_586 (.Y(g7717),.A(g6863),.B(g3206));
NAND2X1 NAND2_587 (.Y(I16467),.A(g10716),.B(g10518));
NAND2X1 NAND2_588 (.Y(I4972),.A(g991),.B(I4971));
NAND2X1 NAND2_589 (.Y(I13554),.A(g8262),.B(I13552));
NAND2X1 NAND2_590 (.Y(I16037),.A(g10427),.B(g2707));
NAND2X1 NAND2_591 (.Y(g8302),.A(I13273),.B(I13274));
NAND2X1 NAND2_592 (.Y(I4943),.A(g324),.B(I4941));
NAND2X1 NAND2_593 (.Y(I5485),.A(g1250),.B(I5484));
NAND2X1 NAND2_594 (.Y(g5527),.A(g3978),.B(g4749));
NAND2X1 NAND2_595 (.Y(I10509),.A(g786),.B(I10507));
NAND2X1 NAND2_596 (.Y(g7599),.A(I12144),.B(I12145));
NAND2X1 NAND2_597 (.Y(I10508),.A(g6221),.B(I10507));
NAND2X1 NAND2_598 (.Y(I6126),.A(g1419),.B(I6124));
NAND2X1 NAND2_599 (.Y(I8671),.A(g814),.B(I8669));
NAND2X1 NAND2_600 (.Y(I6760),.A(g2943),.B(g1448));
NAND2X1 NAND2_601 (.Y(g3626),.A(I6778),.B(I6779));
NAND2X1 NAND2_602 (.Y(I11973),.A(g7001),.B(g1462));
NAND2X1 NAND2_603 (.Y(g2389),.A(I5469),.B(I5470));
NAND2X1 NAND2_604 (.Y(I15617),.A(g10153),.B(I15615));
NAND2X1 NAND2_605 (.Y(g5277),.A(g3734),.B(g4538));
NAND2X1 NAND2_606 (.Y(I5005),.A(g421),.B(g312));
NAND2X1 NAND2_607 (.Y(I6779),.A(g650),.B(I6777));
NAND2X1 NAND2_608 (.Y(I6665),.A(g2792),.B(I6664));
NAND2X1 NAND2_609 (.Y(I8589),.A(g4251),.B(g501));
NAND2X1 NAND2_610 (.Y(g8412),.A(I13545),.B(I13546));
NAND2X1 NAND2_611 (.Y(g2963),.A(I6187),.B(I6188));
NAND2X1 NAND2_612 (.Y(I12045),.A(g6951),.B(g1486));
NAND2X1 NAND2_613 (.Y(I16053),.A(g10371),.B(I16051));
NAND2X1 NAND2_614 (.Y(g2109),.A(I4996),.B(I4997));
NAND2X1 NAND2_615 (.Y(g11418),.A(I17306),.B(I17307));
NAND2X1 NAND2_616 (.Y(I13539),.A(g8157),.B(I13537));
NAND2X1 NAND2_617 (.Y(g10475),.A(I16031),.B(I16032));
NAND2X1 NAND2_618 (.Y(I5324),.A(g1336),.B(I5323));
NAND2X1 NAND2_619 (.Y(I13538),.A(g658),.B(I13537));
NAND2X1 NAND2_620 (.Y(I5469),.A(g1245),.B(I5468));
NAND2X1 NAND2_621 (.Y(I5540),.A(g1023),.B(I5538));
NAND2X1 NAND2_622 (.Y(I17505),.A(g7603),.B(I17503));
NAND2X1 NAND2_623 (.Y(I11241),.A(g6760),.B(g790));
NAND2X1 NAND2_624 (.Y(I8803),.A(g4677),.B(g1113));
NAND2X1 NAND2_625 (.Y(I12061),.A(g6961),.B(I12060));
NAND2X1 NAND2_626 (.Y(I8780),.A(g1137),.B(I8778));
AND2X1 AND_tmp530 (.Y(ttmp530),.A(g6517),.B(g6964));
NAND2X1 NAND_tmp531 (.Y(g8745),.A(g8617),.B(ttmp530));
NAND2X1 NAND2_627 (.Y(I4979),.A(g411),.B(I4978));
NAND2X1 NAND2_628 (.Y(g8109),.A(g5052),.B(g7853));
NAND2X1 NAND2_629 (.Y(g8309),.A(I13308),.B(I13309));
NAND2X1 NAND2_630 (.Y(g6758),.A(I10770),.B(I10771));
NAND2X1 NAND2_631 (.Y(I16009),.A(g2689),.B(I16007));
NAND2X1 NAND2_632 (.Y(I15616),.A(g10043),.B(I15615));
NAND2X1 NAND2_633 (.Y(I8662),.A(g4286),.B(g476));
NAND2X1 NAND2_634 (.Y(I16008),.A(g10424),.B(I16007));
NAND2X1 NAND2_635 (.Y(I13515),.A(g8248),.B(I13513));
NAND2X1 NAND2_636 (.Y(I13991),.A(g622),.B(I13990));
NAND2X1 NAND2_637 (.Y(g11276),.A(I17052),.B(I17053));
NAND2X1 NAND2_638 (.Y(I15900),.A(g10287),.B(I15898));
NAND2X1 NAND2_639 (.Y(g2419),.A(I5501),.B(I5502));
NAND2X1 NAND2_640 (.Y(I16074),.A(g10373),.B(I16072));
NAND2X1 NAND2_641 (.Y(I10769),.A(g5944),.B(g1801));
NAND2X1 NAND2_642 (.Y(I7323),.A(g1231),.B(I7321));
NAND2X1 NAND2_643 (.Y(g7978),.A(g7697),.B(g3038));
NAND2X1 NAND2_644 (.Y(I7875),.A(g4109),.B(g810));
NAND2X1 NAND2_645 (.Y(I8562),.A(g4227),.B(I8561));
NAND2X1 NAND2_646 (.Y(I15892),.A(g10286),.B(I15890));
NAND2X1 NAND2_647 (.Y(g3771),.A(I6989),.B(I6990));
NAND2X1 NAND2_648 (.Y(I8605),.A(g4259),.B(I8604));
NAND2X1 NAND2_649 (.Y(g10153),.A(I15452),.B(I15453));
NAND2X1 NAND2_650 (.Y(g5295),.A(I8762),.B(I8763));
NAND2X1 NAND2_651 (.Y(I8751),.A(g4613),.B(I8750));
NAND2X1 NAND2_652 (.Y(I15907),.A(g6899),.B(I15906));
NAND2X1 NAND2_653 (.Y(I5136),.A(g521),.B(I5135));
NAND2X1 NAND2_654 (.Y(I11263),.A(g826),.B(I11261));
NAND2X1 NAND2_655 (.Y(I14204),.A(g591),.B(I14202));
NAND2X1 NAND2_656 (.Y(g8881),.A(I14210),.B(I14211));
NAND2X1 NAND2_657 (.Y(g2105),.A(I4972),.B(I4973));
AND2X1 AND_tmp532 (.Y(ttmp532),.A(g3071),.B(g3011));
NAND2X1 NAND_tmp533 (.Y(g5557),.A(g4538),.B(ttmp532));
NAND2X1 NAND2_658 (.Y(I5230),.A(g182),.B(I5229));
NAND2X1 NAND2_659 (.Y(I8669),.A(g4831),.B(g814));
NAND2X1 NAND2_660 (.Y(g10474),.A(I16024),.B(I16025));
NAND2X1 NAND2_661 (.Y(I8772),.A(g1133),.B(I8770));
NAND2X1 NAND2_662 (.Y(g2445),.A(I5539),.B(I5540));
NAND2X1 NAND2_663 (.Y(g8006),.A(g5552),.B(g7717));
NAND2X1 NAND2_664 (.Y(I10932),.A(g5555),.B(I10930));
NAND2X1 NAND2_665 (.Y(I17504),.A(g11475),.B(I17503));
NAND2X1 NAND2_666 (.Y(I5137),.A(g525),.B(I5135));
NAND2X1 NAND2_667 (.Y(g8305),.A(I13284),.B(I13285));
NAND2X1 NAND2_668 (.Y(I5891),.A(g750),.B(g2057));
NAND2X1 NAND2_669 (.Y(I13273),.A(g1918),.B(I13272));
NAND2X1 NAND2_670 (.Y(I8480),.A(g4455),.B(I8479));
NAND2X1 NAND2_671 (.Y(g4144),.A(g2160),.B(g3044));
NAND2X1 NAND2_672 (.Y(I15906),.A(g6899),.B(g10302));
NAND2X1 NAND2_673 (.Y(I5342),.A(g315),.B(I5341));
NAND2X1 NAND2_674 (.Y(I13514),.A(g686),.B(I13513));
NAND2X1 NAND2_675 (.Y(g8407),.A(I13522),.B(I13523));
NAND2X1 NAND2_676 (.Y(g4088),.A(I7224),.B(I7225));
NAND2X1 NAND2_677 (.Y(g4488),.A(I7876),.B(I7877));
NAND2X1 NAND2_678 (.Y(g7598),.A(I12137),.B(I12138));
AND2X1 AND_tmp534 (.Y(ttmp534),.A(g1814),.B(g1834));
NAND2X1 NAND_tmp535 (.Y(g3222),.A(g2557),.B(ttmp534));
NAND2X1 NAND2_679 (.Y(I16052),.A(g837),.B(I16051));
NAND2X1 NAND2_680 (.Y(I12127),.A(g7103),.B(I12126));
NAND2X1 NAND2_681 (.Y(g10483),.A(I16087),.B(I16088));
NAND2X1 NAND2_682 (.Y(g8415),.A(I13560),.B(I13561));
NAND2X1 NAND2_683 (.Y(g11415),.A(I17289),.B(I17290));
NAND2X1 NAND2_684 (.Y(g6573),.A(I10508),.B(I10509));
NAND2X1 NAND2_685 (.Y(I5676),.A(g1218),.B(I5675));
NAND2X1 NAND2_686 (.Y(I6778),.A(g2892),.B(I6777));
NAND2X1 NAND2_687 (.Y(g9413),.A(I14613),.B(I14614));
NAND2X1 NAND2_688 (.Y(I8779),.A(g4630),.B(I8778));
NAND2X1 NAND2_689 (.Y(I5592),.A(g1696),.B(I5591));
AND2X1 AND_tmp536 (.Y(ttmp536),.A(g591),.B(g8366));
AND2X1 AND_tmp537 (.Y(ttmp537),.A(g2382),.B(ttmp536));
NAND2X1 NAND_tmp538 (.Y(g8502),.A(g605),.B(ttmp537));
NAND2X1 NAND2_690 (.Y(I15609),.A(g10144),.B(I15607));
NAND2X1 NAND2_691 (.Y(I15608),.A(g10149),.B(I15607));
AND2X1 AND_tmp539 (.Y(ttmp539),.A(g2374),.B(g2382));
NAND2X1 NAND_tmp540 (.Y(g3071),.A(g605),.B(ttmp539));
NAND2X1 NAND2_692 (.Y(g10509),.A(g10436),.B(g6023));
NAND2X1 NAND2_693 (.Y(I17461),.A(g11448),.B(I17459));
NAND2X1 NAND2_694 (.Y(I13506),.A(g8247),.B(I13504));
NAND2X1 NAND2_695 (.Y(I5468),.A(g1245),.B(g999));
NAND2X1 NAND2_696 (.Y(g5219),.A(I8651),.B(I8652));
NAND2X1 NAND2_697 (.Y(I5677),.A(g1223),.B(I5675));
AND2X1 AND_tmp541 (.Y(ttmp541),.A(g8737),.B(g8648));
NAND2X1 NAND_tmp542 (.Y(g8826),.A(g8739),.B(ttmp541));
NAND2X1 NAND2_698 (.Y(I17393),.A(g11415),.B(g11414));
NAND2X1 NAND2_699 (.Y(I5866),.A(g2107),.B(I5865));
NAND2X1 NAND2_700 (.Y(I12126),.A(g7103),.B(g170));
NAND2X1 NAND2_701 (.Y(I4978),.A(g411),.B(g333));
NAND2X1 NAND2_702 (.Y(g7587),.A(I12086),.B(I12087));
NAND2X1 NAND2_703 (.Y(g5286),.A(I8751),.B(I8752));
NAND2X1 NAND2_704 (.Y(g8308),.A(I13301),.B(I13302));
NAND2X1 NAND2_705 (.Y(I7864),.A(g4099),.B(I7863));
NAND2X1 NAND2_706 (.Y(I11981),.A(g6957),.B(I11980));
NAND2X1 NAND2_707 (.Y(I12060),.A(g6961),.B(g1478));
NAND2X1 NAND2_708 (.Y(g5225),.A(I8663),.B(I8664));
NAND2X1 NAND2_709 (.Y(g11538),.A(I17568),.B(I17569));
NAND2X1 NAND2_710 (.Y(I13767),.A(g8417),.B(I13765));
NAND2X1 NAND2_711 (.Y(g10396),.A(I15907),.B(I15908));
NAND2X1 NAND2_712 (.Y(I11262),.A(g6775),.B(I11261));
NAND2X1 NAND2_713 (.Y(I13990),.A(g622),.B(g8688));
NAND2X1 NAND2_714 (.Y(I6224),.A(g2544),.B(g1346));
NAND2X1 NAND2_715 (.Y(I5867),.A(g2105),.B(I5865));
NAND2X1 NAND2_716 (.Y(g2493),.A(g1834),.B(g1840));
NAND2X1 NAND2_717 (.Y(I5893),.A(g2057),.B(I5891));
AND2X1 AND_tmp543 (.Y(ttmp543),.A(g591),.B(g611));
NAND2X1 NAND_tmp544 (.Y(g3062),.A(g2369),.B(ttmp543));
NAND2X1 NAND2_718 (.Y(I13521),.A(g695),.B(g8249));
NAND2X1 NAND2_719 (.Y(I5186),.A(g1515),.B(I5184));
NAND2X1 NAND2_720 (.Y(I6771),.A(g3257),.B(I6770));
NAND2X1 NAND2_721 (.Y(I5325),.A(g1341),.B(I5323));
NAND2X1 NAND2_722 (.Y(I17459),.A(g11449),.B(g11448));
NAND2X1 NAND2_723 (.Y(I9557),.A(g5598),.B(g782));
NAND2X1 NAND2_724 (.Y(g11414),.A(I17282),.B(I17283));
NAND2X1 NAND2_725 (.Y(I12067),.A(g7116),.B(g139));
NAND2X1 NAND2_726 (.Y(I12094),.A(g1490),.B(I12092));
NAND2X1 NAND2_727 (.Y(I4964),.A(g406),.B(g330));
NAND2X1 NAND2_728 (.Y(I13272),.A(g1918),.B(g8158));
NAND2X1 NAND2_729 (.Y(I9948),.A(g1796),.B(I9946));
NAND2X1 NAND2_730 (.Y(g10302),.A(I15717),.B(I15718));
NAND2X1 NAND2_731 (.Y(I16332),.A(g4997),.B(I16330));
NAND2X1 NAND2_732 (.Y(I5106),.A(g435),.B(I5104));
NAND2X1 NAND2_733 (.Y(g8847),.A(g8760),.B(g8683));
NAND2X1 NAND2_734 (.Y(g2257),.A(I5283),.B(I5284));
NAND2X1 NAND2_735 (.Y(I12019),.A(g7119),.B(g166));
NAND2X1 NAND2_736 (.Y(I15441),.A(g10035),.B(g10122));
NAND2X1 NAND2_737 (.Y(I11997),.A(g127),.B(I11995));
NAND2X1 NAND2_738 (.Y(I8739),.A(g4607),.B(I8738));
NAND2X1 NAND2_739 (.Y(I5461),.A(g1003),.B(I5459));
NAND2X1 NAND2_740 (.Y(I13766),.A(g731),.B(I13765));
NAND2X1 NAND2_741 (.Y(I8479),.A(g4455),.B(g3530));
NAND2X1 NAND2_742 (.Y(I17295),.A(g11373),.B(g11369));
NAND2X1 NAND2_743 (.Y(I14271),.A(g8840),.B(I14270));
NAND2X1 NAND2_744 (.Y(I4971),.A(g991),.B(g995));
NAND2X1 NAND2_745 (.Y(g8301),.A(I13266),.B(I13267));
NAND2X1 NAND2_746 (.Y(I6110),.A(g2205),.B(I6109));
NAND2X1 NAND2_747 (.Y(g10482),.A(I16080),.B(I16081));
NAND2X1 NAND2_748 (.Y(g10779),.A(I16468),.B(I16469));
NAND2X1 NAND2_749 (.Y(I6762),.A(g1448),.B(I6760));
NAND2X1 NAND2_750 (.Y(I17289),.A(g11366),.B(I17288));
NAND2X1 NAND2_751 (.Y(I5315),.A(g1032),.B(g1027));
NAND2X1 NAND2_752 (.Y(I17288),.A(g11366),.B(g11363));
NAND2X1 NAND2_753 (.Y(I13859),.A(g1448),.B(I13857));
NAND2X1 NAND2_754 (.Y(g7548),.A(I11981),.B(I11982));
NAND2X1 NAND2_755 (.Y(I13858),.A(g8538),.B(I13857));
NAND2X1 NAND2_756 (.Y(I11996),.A(g7107),.B(I11995));
AND2X1 AND_tmp545 (.Y(ttmp545),.A(g6971),.B(g6964));
NAND2X1 NAND_tmp546 (.Y(g8743),.A(g8617),.B(ttmp545));
NAND2X1 NAND2_757 (.Y(I5880),.A(g2115),.B(I5878));
NAND2X1 NAND2_758 (.Y(g10513),.A(g10441),.B(g5345));
NAND2X1 NAND2_759 (.Y(g8411),.A(I13538),.B(I13539));
NAND2X1 NAND2_760 (.Y(I8626),.A(g511),.B(I8624));
NAND2X1 NAND2_761 (.Y(g10505),.A(g10432),.B(g5938));
NAND2X1 NAND2_762 (.Y(I5612),.A(g1280),.B(I5611));
NAND2X1 NAND2_763 (.Y(g4821),.A(I8179),.B(I8180));
NAND2X1 NAND2_764 (.Y(I12076),.A(g174),.B(I12074));
NAND2X1 NAND2_765 (.Y(I12085),.A(g6980),.B(g1470));
NAND2X1 NAND2_766 (.Y(g7567),.A(I12020),.B(I12021));
NAND2X1 NAND2_767 (.Y(I5128),.A(g1389),.B(I5126));
NAND2X1 NAND2_768 (.Y(I6489),.A(g1227),.B(I6487));
NAND2X1 NAND2_769 (.Y(g7593),.A(I12114),.B(I12115));
NAND2X1 NAND2_770 (.Y(I8778),.A(g4630),.B(g1137));
NAND2X1 NAND2_771 (.Y(g10149),.A(I15442),.B(I15443));
NAND2X1 NAND2_772 (.Y(I13902),.A(g1428),.B(I13900));
NAND2X1 NAND2_773 (.Y(I13301),.A(g1936),.B(I13300));
NAND2X1 NAND2_774 (.Y(g3215),.A(g2564),.B(g1822));
AND2X1 AND_tmp547 (.Y(ttmp547),.A(g7562),.B(g6974));
AND2X1 AND_tmp548 (.Y(ttmp548),.A(g7011),.B(ttmp547));
NAND2X1 NAND_tmp549 (.Y(g7996),.A(g7574),.B(ttmp548));
NAND2X1 NAND2_775 (.Y(I4985),.A(g999),.B(g1003));
NAND2X1 NAND2_776 (.Y(I14444),.A(g1834),.B(I14442));
AND2X1 AND_tmp550 (.Y(ttmp550),.A(g7562),.B(g7550));
AND2X1 AND_tmp551 (.Y(ttmp551),.A(g7011),.B(ttmp550));
NAND2X1 NAND_tmp552 (.Y(g8000),.A(g7574),.B(ttmp551));
NAND2X1 NAND2_777 (.Y(I5166),.A(g1499),.B(I5164));
NAND2X1 NAND2_778 (.Y(I17460),.A(g11449),.B(I17459));
NAND2X1 NAND2_779 (.Y(g3008),.A(g2444),.B(g878));
NAND2X1 NAND2_780 (.Y(I6836),.A(g3287),.B(g806));
NAND2X1 NAND2_781 (.Y(I5529),.A(g1265),.B(I5528));
NAND2X1 NAND2_782 (.Y(g10229),.A(I15608),.B(I15609));
NAND2X1 NAND2_783 (.Y(I13661),.A(g8322),.B(I13659));
NAND2X1 NAND2_784 (.Y(I13895),.A(g1436),.B(I13893));
NAND2X1 NAND2_785 (.Y(g2303),.A(I5342),.B(I5343));
NAND2X1 NAND2_786 (.Y(I12039),.A(g6990),.B(I12038));
NAND2X1 NAND2_787 (.Y(g5592),.A(I9007),.B(I9008));
NAND2X1 NAND2_788 (.Y(I12038),.A(g6990),.B(g1466));
NAND2X1 NAND2_789 (.Y(g3322),.A(I6488),.B(I6489));
NAND2X1 NAND2_790 (.Y(I8561),.A(g4227),.B(g491));
NAND2X1 NAND2_791 (.Y(I8527),.A(g4879),.B(g481));
NAND2X1 NAND2_792 (.Y(I12143),.A(g7089),.B(g158));
NAND2X1 NAND2_793 (.Y(I5619),.A(g1766),.B(I5618));
NAND2X1 NAND2_794 (.Y(g10386),.A(I15879),.B(I15880));
NAND2X1 NAND2_795 (.Y(I11980),.A(g6957),.B(g1482));
NAND2X1 NAND2_796 (.Y(I6837),.A(g3287),.B(I6836));
NAND2X1 NAND2_797 (.Y(I4973),.A(g995),.B(I4971));
NAND2X1 NAND2_798 (.Y(I13888),.A(g1440),.B(I13886));
NAND2X1 NAND2_799 (.Y(g7558),.A(I12003),.B(I12004));
NAND2X1 NAND2_800 (.Y(I17494),.A(g3623),.B(I17492));
NAND2X1 NAND2_801 (.Y(g11491),.A(I17493),.B(I17494));
NAND2X1 NAND2_802 (.Y(I16045),.A(g833),.B(I16044));
NAND2X1 NAND2_803 (.Y(I7684),.A(g1023),.B(I7683));
NAND2X1 NAND2_804 (.Y(g4130),.A(g3044),.B(g2518));
NAND2X1 NAND2_805 (.Y(I8771),.A(g4619),.B(I8770));
NAND2X1 NAND2_806 (.Y(I13546),.A(g8259),.B(I13544));
NAND2X1 NAND2_807 (.Y(I13089),.A(g8006),.B(g1840));
NAND2X1 NAND2_808 (.Y(g2117),.A(I5024),.B(I5025));
NAND2X1 NAND2_809 (.Y(g5119),.A(I8514),.B(I8515));
NAND2X1 NAND2_810 (.Y(g5319),.A(I8804),.B(I8805));
NAND2X1 NAND2_811 (.Y(I15899),.A(g857),.B(I15898));
NAND2X1 NAND2_812 (.Y(I5606),.A(g1153),.B(I5604));
NAND2X1 NAND2_813 (.Y(I15898),.A(g857),.B(g10287));
NAND2X1 NAND2_814 (.Y(I16032),.A(g10368),.B(I16030));
NAND2X1 NAND2_815 (.Y(I17401),.A(g11418),.B(I17400));
NAND2X1 NAND2_816 (.Y(I13659),.A(g1945),.B(g8322));
NAND2X1 NAND2_817 (.Y(I8738),.A(g4607),.B(g1121));
NAND2X1 NAND2_818 (.Y(I13250),.A(g8148),.B(I13248));
NAND2X1 NAND2_819 (.Y(I15718),.A(g10229),.B(I15716));
NAND2X1 NAND2_820 (.Y(I9008),.A(g1791),.B(I9006));
NAND2X1 NAND2_821 (.Y(I6176),.A(g2177),.B(g197));
NAND2X1 NAND2_822 (.Y(I7865),.A(g774),.B(I7863));
NAND2X1 NAND2_823 (.Y(g5274),.A(I8729),.B(I8730));
NAND2X1 NAND2_824 (.Y(I5341),.A(g315),.B(g426));
NAND2X1 NAND2_825 (.Y(I17305),.A(g11381),.B(g11377));
NAND2X1 NAND2_826 (.Y(I17053),.A(g11249),.B(I17051));
NAND2X1 NAND2_827 (.Y(g5125),.A(I8528),.B(I8529));
NAND2X1 NAND2_828 (.Y(I12216),.A(g2518),.B(I12214));
NAND2X1 NAND2_829 (.Y(I6225),.A(g2544),.B(I6224));
NAND2X1 NAND2_830 (.Y(I5879),.A(g2120),.B(I5878));
NAND2X1 NAND2_831 (.Y(g3221),.A(g1834),.B(g2564));
NAND2X1 NAND2_832 (.Y(I14270),.A(g8840),.B(g1822));
NAND2X1 NAND2_833 (.Y(I6124),.A(g2215),.B(g1419));
NAND2X1 NAND2_834 (.Y(I6324),.A(g1864),.B(I6322));
NAND2X1 NAND2_835 (.Y(I13867),.A(g8523),.B(g1403));
NAND2X1 NAND2_836 (.Y(I13894),.A(g8529),.B(I13893));
NAND2X1 NAND2_837 (.Y(I6469),.A(g2479),.B(I6467));
NAND2X1 NAND2_838 (.Y(I8663),.A(g4286),.B(I8662));
NAND2X1 NAND2_839 (.Y(g7523),.A(I11908),.B(I11909));
NAND2X1 NAND2_840 (.Y(I6177),.A(g2177),.B(I6176));
NAND2X1 NAND2_841 (.Y(g5187),.A(I8590),.B(I8591));
NAND2X1 NAND2_842 (.Y(I6287),.A(g2091),.B(g981));
NAND2X1 NAND2_843 (.Y(I8762),.A(g4616),.B(I8761));
NAND2X1 NAND2_844 (.Y(I15871),.A(g10358),.B(I15870));
AND2X1 AND_tmp553 (.Y(ttmp553),.A(g8541),.B(g8760));
NAND2X1 NAND_tmp554 (.Y(g8840),.A(g8542),.B(ttmp553));
NAND2X1 NAND2_845 (.Y(g2250),.A(I5264),.B(I5265));
NAND2X1 NAND2_846 (.Y(I8590),.A(g4251),.B(I8589));
NAND2X1 NAND2_847 (.Y(I6199),.A(g2525),.B(g766));
NAND2X1 NAND2_848 (.Y(I14218),.A(g605),.B(I14216));
NAND2X1 NAND2_849 (.Y(g8190),.A(g6027),.B(g7978));
NAND2X1 NAND2_850 (.Y(I5284),.A(g762),.B(I5282));
NAND2X1 NAND2_851 (.Y(I17485),.A(g11384),.B(g11474));
NAND2X1 NAND2_852 (.Y(I4965),.A(g406),.B(I4964));
NAND2X1 NAND2_853 (.Y(I5591),.A(g1696),.B(g1703));
NAND2X1 NAND2_854 (.Y(g8501),.A(g3760),.B(g8366));
NAND2X1 NAND2_855 (.Y(I15451),.A(g10058),.B(g10051));
NAND2X1 NAND2_856 (.Y(g8942),.A(g8823),.B(g4921));
NAND2X1 NAND2_857 (.Y(I13877),.A(g8535),.B(I13876));
NAND2X1 NAND2_858 (.Y(g7269),.A(I11509),.B(I11510));
NAND2X1 NAND2_859 (.Y(I4996),.A(g416),.B(I4995));
NAND2X1 NAND2_860 (.Y(I6144),.A(g1976),.B(I6143));
NAND2X1 NAND2_861 (.Y(I17567),.A(g11496),.B(g1610));
NAND2X1 NAND2_862 (.Y(g7572),.A(I12039),.B(I12040));
NAND2X1 NAND2_863 (.Y(I6207),.A(g2534),.B(g802));
NAND2X1 NAND2_864 (.Y(I14277),.A(g8847),.B(g1828));
NAND2X1 NAND2_865 (.Y(I16059),.A(g841),.B(I16058));
NAND2X1 NAND2_866 (.Y(I16025),.A(g2701),.B(I16023));
NAND2X1 NAND2_867 (.Y(I8563),.A(g491),.B(I8561));
NAND2X1 NAND2_868 (.Y(g3524),.A(g3209),.B(g3221));
NAND2X1 NAND2_869 (.Y(I16058),.A(g841),.B(g10372));
NAND2X1 NAND2_870 (.Y(I5204),.A(g374),.B(I5202));
NAND2X1 NAND2_871 (.Y(I6488),.A(g2306),.B(I6487));
AND2X1 AND_tmp555 (.Y(ttmp555),.A(g2310),.B(g3003));
AND2X1 AND_tmp556 (.Y(ttmp556),.A(g3056),.B(ttmp555));
NAND2X1 NAND_tmp557 (.Y(g3818),.A(g3071),.B(ttmp556));
NAND2X1 NAND2_872 (.Y(I16044),.A(g833),.B(g10370));
NAND2X1 NAND2_873 (.Y(g3717),.A(I6880),.B(I6881));
NAND2X1 NAND2_874 (.Y(I13077),.A(g1872),.B(I13076));
NAND2X1 NAND2_875 (.Y(g10043),.A(I15257),.B(I15258));
NAND2X1 NAND2_876 (.Y(I11280),.A(g6485),.B(I11278));
NAND2X1 NAND2_877 (.Y(I6825),.A(g3281),.B(g770));
NAND2X1 NAND2_878 (.Y(I4997),.A(g309),.B(I4995));
NAND2X1 NAND2_879 (.Y(I13300),.A(g1936),.B(g8162));
NAND2X1 NAND2_880 (.Y(I5323),.A(g1336),.B(g1341));
NAND2X1 NAND2_881 (.Y(I6136),.A(g2496),.B(g378));
NAND2X1 NAND2_882 (.Y(g5935),.A(I9558),.B(I9559));
NAND2X1 NAND2_883 (.Y(I5528),.A(g1265),.B(g1015));
NAND2X1 NAND2_884 (.Y(I6806),.A(g3268),.B(I6805));
NAND2X1 NAND2_885 (.Y(I5530),.A(g1015),.B(I5528));
NAND2X1 NAND2_886 (.Y(g10886),.A(g10807),.B(g10805));
NAND2X1 NAND2_887 (.Y(g3106),.A(I6323),.B(I6324));
NAND2X1 NAND2_888 (.Y(I13876),.A(g8535),.B(g1444));
NAND2X1 NAND2_889 (.Y(I6322),.A(g2050),.B(g1864));
NAND2X1 NAND2_890 (.Y(g3061),.A(g611),.B(g2374));
NAND2X1 NAND2_891 (.Y(g2439),.A(g1814),.B(g1828));
AND2X1 AND_tmp558 (.Y(ttmp558),.A(g7279),.B(g7369));
AND2X1 AND_tmp559 (.Y(ttmp559),.A(g7395),.B(ttmp558));
NAND2X1 NAND_tmp560 (.Y(g7947),.A(g7390),.B(ttmp559));
NAND2X1 NAND2_892 (.Y(I9576),.A(g818),.B(I9574));
NAND2X1 NAND2_893 (.Y(I13660),.A(g1945),.B(I13659));
NAND2X1 NAND2_894 (.Y(g3200),.A(g1822),.B(g2061));
NAND2X1 NAND2_895 (.Y(g4374),.A(I7684),.B(I7685));
NAND2X1 NAND2_896 (.Y(I11916),.A(g1494),.B(I11914));
NAND2X1 NAND2_897 (.Y(I5372),.A(g971),.B(I5371));
NAND2X1 NAND2_898 (.Y(g3003),.A(g599),.B(g2399));
NAND2X1 NAND2_899 (.Y(g8627),.A(I13887),.B(I13888));
NAND2X1 NAND2_900 (.Y(I5618),.A(g1766),.B(g1771));
NAND2X1 NAND2_901 (.Y(I6137),.A(g2496),.B(I6136));
NAND2X1 NAND2_902 (.Y(I5343),.A(g426),.B(I5341));
NAND2X1 NAND2_903 (.Y(I5282),.A(g758),.B(g762));
NAND2X1 NAND2_904 (.Y(I13307),.A(g8190),.B(g617));
NAND2X1 NAND2_905 (.Y(I13076),.A(g1872),.B(g7963));
NAND2X1 NAND2_906 (.Y(I6807),.A(g471),.B(I6805));
NAND2X1 NAND2_907 (.Y(I11243),.A(g790),.B(I11241));
NAND2X1 NAND2_908 (.Y(I17585),.A(g11354),.B(I17584));
NAND2X1 NAND2_909 (.Y(I12137),.A(g7110),.B(I12136));
NAND2X1 NAND2_910 (.Y(I7564),.A(g654),.B(I7562));
NAND2X1 NAND2_911 (.Y(g2970),.A(I6200),.B(I6201));
NAND2X1 NAND2_912 (.Y(g10144),.A(I15431),.B(I15432));
NAND2X1 NAND2_913 (.Y(I8788),.A(g1141),.B(I8786));
NAND2X1 NAND2_914 (.Y(g7054),.A(I11242),.B(I11243));
NAND2X1 NAND2_915 (.Y(I17052),.A(g10923),.B(I17051));
NAND2X1 NAND2_916 (.Y(g2120),.A(I5035),.B(I5036));
NAND2X1 NAND2_917 (.Y(g8616),.A(I13868),.B(I13869));
NAND2X1 NAND2_918 (.Y(I5202),.A(g369),.B(g374));
NAND2X1 NAND2_919 (.Y(I16088),.A(g10375),.B(I16086));
NAND2X1 NAND2_920 (.Y(I16024),.A(g10426),.B(I16023));
NAND2X1 NAND2_921 (.Y(g11490),.A(I17486),.B(I17487));
NAND2X1 NAND2_922 (.Y(I5518),.A(g1019),.B(I5516));
AND2X1 AND_tmp561 (.Y(ttmp561),.A(g4806),.B(g4073));
NAND2X1 NAND_tmp562 (.Y(g5118),.A(g2439),.B(ttmp561));
NAND2X1 NAND2_923 (.Y(I12021),.A(g166),.B(I12019));
NOR2X1 NOR2_0 (.Y(g6392),.A(g5859),.B(g5938));
NOR2X1 NOR2_1 (.Y(g5938),.A(g2764),.B(g4988));
NOR2X1 NOR2_2 (.Y(g2478),.A(g1610),.B(g1737));
NOR2X1 NOR2_3 (.Y(g10374),.A(g10347),.B(g3463));
OR2X1 OR_tmp563 (.Y(ttmp563),.A(g2586),.B(g3776));
OR2X1 OR_tmp564 (.Y(ttmp564),.A(g3800),.B(ttmp563));
NOR2X1 NOR_tmp565 (.Y(g4278),.A(g2593),.B(ttmp564));
NOR2X1 NOR2_4 (.Y(g10424),.A(g10292),.B(g4620));
NOR2X1 NOR2_5 (.Y(g10383),.A(g10318),.B(g2998));
NOR2X1 NOR2_6 (.Y(g3118),.A(g2521),.B(g2514));
NOR2X1 NOR2_7 (.Y(g9815),.A(g9392),.B(g9367));
NOR2X1 NOR2_8 (.Y(g11077),.A(g10970),.B(g10971));
OR2X1 OR_tmp566 (.Y(ttmp566),.A(g9274),.B(g9292));
NOR2X1 NOR_tmp567 (.Y(g9746),.A(g9454),.B(ttmp566));
OR2X1 OR_tmp568 (.Y(ttmp568),.A(g2354),.B(g2353));
NOR2X1 NOR_tmp569 (.Y(g3879),.A(g3141),.B(ttmp568));
NOR2X1 NOR2_9 (.Y(g10285),.A(g10276),.B(g3566));
NOR2X1 NOR2_10 (.Y(g11480),.A(g11456),.B(g4567));
NOR2X1 NOR2_11 (.Y(g4076),.A(g1707),.B(g2864));
NOR2X1 NOR2_12 (.Y(g10570),.A(g10542),.B(g10324));
NOR2X1 NOR2_13 (.Y(g10239),.A(g9317),.B(g10179));
NOR2X1 NOR2_14 (.Y(g10594),.A(g10480),.B(g10521));
NOR2X1 NOR2_15 (.Y(g9426),.A(g9052),.B(g9030));
NOR2X1 NOR2_16 (.Y(g10382),.A(g10314),.B(g2998));
OR2X1 OR_tmp570 (.Y(ttmp570),.A(g2662),.B(g3479));
OR2X1 OR_tmp571 (.Y(ttmp571),.A(g3501),.B(ttmp570));
NOR2X1 NOR_tmp572 (.Y(g4672),.A(g2669),.B(ttmp571));
NOR2X1 NOR2_17 (.Y(g5360),.A(g2071),.B(g4225));
OR2X1 OR_tmp573 (.Y(ttmp573),.A(g9223),.B(I14596));
OR2X1 OR_tmp574 (.Y(ttmp574),.A(g9010),.B(ttmp573));
NOR2X1 NOR_tmp575 (.Y(g9387),.A(g9240),.B(ttmp574));
NOR2X1 NOR2_18 (.Y(g10438),.A(g10356),.B(g3566));
OR2X1 OR_tmp576 (.Y(ttmp576),.A(g2662),.B(g2655));
OR2X1 OR_tmp577 (.Y(ttmp577),.A(g3077),.B(ttmp576));
NOR2X1 NOR_tmp578 (.Y(g4613),.A(g3491),.B(ttmp577));
OR2X1 OR_tmp579 (.Y(ttmp579),.A(g9223),.B(I14602));
OR2X1 OR_tmp580 (.Y(ttmp580),.A(g9010),.B(ttmp579));
NOR2X1 NOR_tmp581 (.Y(g9391),.A(g9240),.B(ttmp580));
OR2X1 OR_tmp582 (.Y(ttmp582),.A(g3408),.B(g3628));
NOR2X1 NOR_tmp583 (.Y(g4572),.A(g3419),.B(ttmp582));
OR2X1 OR_tmp584 (.Y(ttmp584),.A(g9274),.B(g9292));
NOR2X1 NOR_tmp585 (.Y(g9757),.A(g9454),.B(ttmp584));
NOR2X1 NOR2_19 (.Y(g9416),.A(g9052),.B(g9030));
OR2X1 OR_tmp586 (.Y(ttmp586),.A(g9579),.B(I15033));
OR2X1 OR_tmp587 (.Y(ttmp587),.A(g9519),.B(ttmp586));
NOR2X1 NOR_tmp588 (.Y(g9874),.A(g9536),.B(ttmp587));
NOR2X1 NOR2_20 (.Y(g9654),.A(g9125),.B(g9173));
OR2X1 OR_tmp589 (.Y(ttmp589),.A(g9557),.B(I15051));
OR2X1 OR_tmp590 (.Y(ttmp590),.A(g9751),.B(ttmp589));
NOR2X1 NOR_tmp591 (.Y(g9880),.A(g9536),.B(ttmp590));
OR2X1 OR_tmp592 (.Y(ttmp592),.A(g2586),.B(g3776));
OR2X1 OR_tmp593 (.Y(ttmp593),.A(g3292),.B(ttmp592));
NOR2X1 NOR_tmp594 (.Y(g4873),.A(g2593),.B(ttmp593));
NOR2X1 NOR2_21 (.Y(g2807),.A(g22),.B(g2320));
NOR2X1 NOR2_22 (.Y(g10441),.A(g10351),.B(g3566));
OR2X1 OR_tmp595 (.Y(ttmp595),.A(g2662),.B(g2655));
OR2X1 OR_tmp596 (.Y(ttmp596),.A(g3501),.B(ttmp595));
NOR2X1 NOR_tmp597 (.Y(g4639),.A(g2669),.B(ttmp596));
NOR2X1 NOR2_23 (.Y(g10435),.A(g10332),.B(g3507));
NOR2X1 NOR2_24 (.Y(g10849),.A(g10739),.B(g3903));
OR2X1 OR_tmp598 (.Y(ttmp598),.A(g9173),.B(g9151));
OR2X1 OR_tmp599 (.Y(ttmp599),.A(g9125),.B(ttmp598));
NOR2X1 NOR_tmp600 (.Y(g9606),.A(g9111),.B(ttmp599));
OR2X1 OR_tmp601 (.Y(ttmp601),.A(g9566),.B(I15048));
OR2X1 OR_tmp602 (.Y(ttmp602),.A(g9747),.B(ttmp601));
NOR2X1 NOR_tmp603 (.Y(g9879),.A(g9536),.B(ttmp602));
NOR2X1 NOR2_25 (.Y(g9506),.A(g9052),.B(g9030));
NOR2X1 NOR2_26 (.Y(g6155),.A(g4974),.B(g2864));
NOR2X1 NOR2_27 (.Y(g6355),.A(g6032),.B(g6023));
NOR2X1 NOR2_28 (.Y(g9615),.A(g9052),.B(g9030));
NOR2X1 NOR2_29 (.Y(g10371),.A(g10344),.B(g3463));
NOR2X1 NOR2_30 (.Y(g9591),.A(g9125),.B(g9151));
NOR2X1 NOR2_31 (.Y(g10359),.A(g10227),.B(g4620));
NOR2X1 NOR2_32 (.Y(g10434),.A(g10352),.B(g3566));
NOR2X1 NOR2_33 (.Y(g10358),.A(g10226),.B(g4620));
OR2X1 OR_tmp604 (.Y(ttmp604),.A(g9274),.B(g9292));
NOR2X1 NOR_tmp605 (.Y(g9750),.A(g9454),.B(ttmp604));
NOR2X1 NOR2_34 (.Y(g10291),.A(g10247),.B(g3113));
OR2X1 OR_tmp606 (.Y(ttmp606),.A(g2586),.B(g2579));
OR2X1 OR_tmp607 (.Y(ttmp607),.A(g3292),.B(ttmp606));
NOR2X1 NOR_tmp608 (.Y(g4227),.A(g3793),.B(ttmp607));
OR2X1 OR_tmp609 (.Y(ttmp609),.A(g9223),.B(I14776));
OR2X1 OR_tmp610 (.Y(ttmp610),.A(g9010),.B(ttmp609));
NOR2X1 NOR_tmp611 (.Y(g9655),.A(g9240),.B(ttmp610));
OR2X1 OR_tmp612 (.Y(ttmp612),.A(g9223),.B(I14607));
OR2X1 OR_tmp613 (.Y(ttmp613),.A(g9010),.B(ttmp612));
NOR2X1 NOR_tmp614 (.Y(g9410),.A(g9240),.B(ttmp613));
OR2X1 OR_tmp615 (.Y(ttmp615),.A(g9173),.B(g9151));
OR2X1 OR_tmp616 (.Y(ttmp616),.A(g9125),.B(ttmp615));
NOR2X1 NOR_tmp617 (.Y(g9667),.A(g9111),.B(ttmp616));
NOR2X1 NOR2_35 (.Y(g10563),.A(g10539),.B(g10322));
NOR2X1 NOR2_36 (.Y(g9776),.A(g9392),.B(g9367));
NOR2X1 NOR2_37 (.Y(g10324),.A(g9317),.B(g10244));
OR2X1 OR_tmp618 (.Y(ttmp618),.A(g3419),.B(g3408));
NOR2X1 NOR_tmp619 (.Y(g4455),.A(g3543),.B(ttmp618));
OR2X1 OR_tmp620 (.Y(ttmp620),.A(g9560),.B(I15045));
OR2X1 OR_tmp621 (.Y(ttmp621),.A(g9754),.B(ttmp620));
NOR2X1 NOR_tmp622 (.Y(g9878),.A(g9536),.B(ttmp621));
NOR2X1 NOR2_38 (.Y(g10360),.A(g10277),.B(g3566));
OR2X1 OR_tmp623 (.Y(ttmp623),.A(g9563),.B(I15057));
OR2X1 OR_tmp624 (.Y(ttmp624),.A(g9742),.B(ttmp623));
NOR2X1 NOR_tmp625 (.Y(g9882),.A(g9536),.B(ttmp624));
NOR2X1 NOR2_39 (.Y(g10370),.A(g10343),.B(g3463));
OR2X1 OR_tmp626 (.Y(ttmp626),.A(g3485),.B(g2655));
OR2X1 OR_tmp627 (.Y(ttmp627),.A(g3077),.B(ttmp626));
NOR2X1 NOR_tmp628 (.Y(g4605),.A(g2669),.B(ttmp627));
NOR2X1 NOR2_40 (.Y(g10420),.A(g10329),.B(g3744));
NOR2X1 NOR2_41 (.Y(g10562),.A(g10483),.B(g10529));
NOR2X1 NOR2_42 (.Y(g10427),.A(g10296),.B(g4620));
NOR2X1 NOR2_43 (.Y(g5780),.A(g2112),.B(g4921));
NOR2X1 NOR2_44 (.Y(g10385),.A(g10321),.B(g2998));
NOR2X1 NOR2_45 (.Y(g10376),.A(g10323),.B(g3113));
NOR2X1 NOR2_46 (.Y(g10426),.A(g10294),.B(g4620));
OR2X1 OR_tmp629 (.Y(ttmp629),.A(g2662),.B(g3479));
OR2X1 OR_tmp630 (.Y(ttmp630),.A(g3077),.B(ttmp629));
NOR2X1 NOR_tmp631 (.Y(g4601),.A(g2669),.B(ttmp630));
NOR2X1 NOR2_47 (.Y(g5573),.A(g4117),.B(g4432));
NOR2X1 NOR2_48 (.Y(g9808),.A(g9392),.B(g9367));
NOR2X1 NOR2_49 (.Y(g5999),.A(g2753),.B(g4953));
OR2X1 OR_tmp632 (.Y(ttmp632),.A(g9274),.B(g9292));
NOR2X1 NOR_tmp633 (.Y(g9759),.A(g9454),.B(ttmp632));
NOR2X1 NOR2_50 (.Y(g6037),.A(g3305),.B(g5614));
NOR2X1 NOR2_51 (.Y(g10287),.A(g10275),.B(g3463));
NOR2X1 NOR2_52 (.Y(g5034),.A(g3524),.B(g4593));
OR2X1 OR_tmp634 (.Y(ttmp634),.A(g9223),.B(I14585));
OR2X1 OR_tmp635 (.Y(ttmp635),.A(g9010),.B(ttmp634));
NOR2X1 NOR_tmp636 (.Y(g9362),.A(g9240),.B(ttmp635));
OR2X1 OR_tmp637 (.Y(ttmp637),.A(g9573),.B(I15054));
OR2X1 OR_tmp638 (.Y(ttmp638),.A(g9516),.B(ttmp637));
NOR2X1 NOR_tmp639 (.Y(g9881),.A(g9536),.B(ttmp638));
NOR2X1 NOR2_53 (.Y(g10443),.A(g10353),.B(g3566));
NOR2X1 NOR2_54 (.Y(g10286),.A(g10271),.B(g3463));
OR2X1 OR_tmp640 (.Y(ttmp640),.A(g3261),.B(g2500));
NOR2X1 NOR_tmp641 (.Y(g4276),.A(g4065),.B(ttmp640));
OR2X1 OR_tmp642 (.Y(ttmp642),.A(g2662),.B(g3479));
OR2X1 OR_tmp643 (.Y(ttmp643),.A(g3077),.B(ttmp642));
NOR2X1 NOR_tmp644 (.Y(g4616),.A(g3491),.B(ttmp643));
NOR2X1 NOR2_55 (.Y(g10363),.A(g10355),.B(g3566));
NOR2X1 NOR2_56 (.Y(g2862),.A(g2315),.B(g2305));
NOR2X1 NOR2_57 (.Y(g10373),.A(g10346),.B(g3463));
NOR2X1 NOR2_58 (.Y(g10423),.A(g10290),.B(g4620));
OR2X1 OR_tmp645 (.Y(ttmp645),.A(g9274),.B(g9292));
NOR2X1 NOR_tmp646 (.Y(g9758),.A(g9454),.B(ttmp645));
OR2X1 OR_tmp647 (.Y(ttmp647),.A(g9173),.B(g9151));
NOR2X1 NOR_tmp648 (.Y(g9589),.A(g9125),.B(ttmp647));
NOR2X1 NOR2_59 (.Y(g9803),.A(g9392),.B(g9367));
NOR2X1 NOR2_60 (.Y(g10430),.A(g10349),.B(g3566));
NOR2X1 NOR2_61 (.Y(g9421),.A(g9052),.B(g9030));
NOR2X1 NOR2_62 (.Y(g10362),.A(g10228),.B(g3507));
NOR2X1 NOR2_63 (.Y(g2791),.A(g2187),.B(g750));
NOR2X1 NOR2_64 (.Y(g9817),.A(g9392),.B(g9367));
OR2X1 OR_tmp649 (.Y(ttmp649),.A(g9173),.B(g9151));
OR2X1 OR_tmp650 (.Y(ttmp650),.A(g9125),.B(ttmp649));
NOR2X1 NOR_tmp651 (.Y(g9605),.A(g9111),.B(ttmp650));
NOR2X1 NOR2_65 (.Y(g10372),.A(g10345),.B(g3463));
NOR2X1 NOR2_66 (.Y(g9669),.A(g9392),.B(g9367));
NOR2X1 NOR2_67 (.Y(g10422),.A(g10289),.B(g4620));
NOR2X1 NOR2_68 (.Y(g10436),.A(g10354),.B(g3566));
OR2X1 OR_tmp652 (.Y(ttmp652),.A(g2299),.B(g2031));
OR2X1 OR_tmp653 (.Y(ttmp653),.A(g4787),.B(ttmp652));
NOR2X1 NOR_tmp654 (.Y(g5556),.A(g2695),.B(ttmp653));
OR2X1 OR_tmp655 (.Y(ttmp655),.A(g3784),.B(g2579));
OR2X1 OR_tmp656 (.Y(ttmp656),.A(g3800),.B(ttmp655));
NOR2X1 NOR_tmp657 (.Y(g4286),.A(g2593),.B(ttmp656));
NOR2X1 NOR2_69 (.Y(g4974),.A(g4502),.B(g3714));
NOR2X1 NOR2_70 (.Y(g9779),.A(g9392),.B(g9367));
NOR2X1 NOR2_71 (.Y(g9423),.A(g9052),.B(g9030));
NOR2X1 NOR2_72 (.Y(g5350),.A(g4163),.B(g4872));
OR2X1 OR_tmp658 (.Y(ttmp658),.A(g9223),.B(I14582));
OR2X1 OR_tmp659 (.Y(ttmp659),.A(g9010),.B(ttmp658));
NOR2X1 NOR_tmp660 (.Y(g9361),.A(g9240),.B(ttmp659));
OR2X1 OR_tmp661 (.Y(ttmp661),.A(g1651),.B(g1648));
OR2X1 OR_tmp662 (.Y(ttmp662),.A(g1645),.B(ttmp661));
NOR2X1 NOR_tmp663 (.Y(g2459),.A(g1642),.B(ttmp662));
NOR2X1 NOR2_73 (.Y(g10381),.A(g10310),.B(g2998));
OR2X1 OR_tmp664 (.Y(ttmp664),.A(g3784),.B(g3776));
OR2X1 OR_tmp665 (.Y(ttmp665),.A(g3292),.B(ttmp664));
NOR2X1 NOR_tmp666 (.Y(g4259),.A(g3793),.B(ttmp665));
NOR2X1 NOR2_74 (.Y(g10522),.A(g10486),.B(g10239));
NOR2X1 NOR2_75 (.Y(g5392),.A(g3369),.B(g4258));
OR2X1 OR_tmp667 (.Y(ttmp667),.A(g2410),.B(g2538));
NOR2X1 NOR_tmp668 (.Y(g4122),.A(g3291),.B(ttmp667));
NOR2X1 NOR2_76 (.Y(g6023),.A(g2763),.B(g4975));
NOR2X1 NOR2_77 (.Y(g3462),.A(g2187),.B(g2795));
OR2X1 OR_tmp669 (.Y(ttmp669),.A(g3784),.B(g3776));
OR2X1 OR_tmp670 (.Y(ttmp670),.A(g3292),.B(ttmp669));
NOR2X1 NOR_tmp671 (.Y(g4218),.A(g2593),.B(ttmp670));
OR2X1 OR_tmp672 (.Y(ttmp672),.A(g2586),.B(g2579));
OR2X1 OR_tmp673 (.Y(ttmp673),.A(g3800),.B(ttmp672));
NOR2X1 NOR_tmp674 (.Y(g4267),.A(g2593),.B(ttmp673));
OR2X1 OR_tmp675 (.Y(ttmp675),.A(g3485),.B(g2655));
OR2X1 OR_tmp676 (.Y(ttmp676),.A(g3501),.B(ttmp675));
NOR2X1 NOR_tmp677 (.Y(g4677),.A(g2669),.B(ttmp676));
NOR2X1 NOR2_78 (.Y(g9646),.A(g9125),.B(g9151));
NOR2X1 NOR2_79 (.Y(g2863),.A(g2316),.B(g2309));
OR2X1 OR_tmp678 (.Y(ttmp678),.A(g9223),.B(I14751));
OR2X1 OR_tmp679 (.Y(ttmp679),.A(g9010),.B(ttmp678));
NOR2X1 NOR_tmp680 (.Y(g9616),.A(g9240),.B(ttmp679));
NOR2X1 NOR2_80 (.Y(g6032),.A(g3430),.B(g5039));
OR2X1 OR_tmp681 (.Y(ttmp681),.A(g9173),.B(g9151));
OR2X1 OR_tmp682 (.Y(ttmp682),.A(g9125),.B(ttmp681));
NOR2X1 NOR_tmp683 (.Y(g9647),.A(g9111),.B(ttmp682));
NOR2X1 NOR2_81 (.Y(g5859),.A(g3362),.B(g4943));
NOR2X1 NOR2_82 (.Y(g10433),.A(g10330),.B(g3507));
NOR2X1 NOR2_83 (.Y(g10368),.A(g10342),.B(g3463));
OR2X1 OR_tmp684 (.Y(ttmp684),.A(g3784),.B(g2579));
OR2X1 OR_tmp685 (.Y(ttmp685),.A(g3292),.B(ttmp684));
NOR2X1 NOR_tmp686 (.Y(g4251),.A(g3793),.B(ttmp685));
OR2X1 OR_tmp687 (.Y(ttmp687),.A(g9576),.B(I15039));
OR2X1 OR_tmp688 (.Y(ttmp688),.A(g9522),.B(ttmp687));
NOR2X1 NOR_tmp689 (.Y(g9876),.A(g9536),.B(ttmp688));
OR2X1 OR_tmp690 (.Y(ttmp690),.A(g9223),.B(I14779));
OR2X1 OR_tmp691 (.Y(ttmp691),.A(g9010),.B(ttmp690));
NOR2X1 NOR_tmp692 (.Y(g9656),.A(g9240),.B(ttmp691));
NOR2X1 NOR2_84 (.Y(g8303),.A(g8209),.B(g4811));
NOR2X1 NOR2_85 (.Y(g10429),.A(g10326),.B(g3507));
OR2X1 NOR2_86 (.Y(g10428),.A(g10335),.B(g4620));
NOR2X1 OR_tmp693 (.Y(ttmp693),.A(g2586),.B(g3776));
OR2X1 OR_tmp694 (.Y(ttmp694),.A(g3292),.B(ttmp693));
NOR2X1 NOR_tmp695 (.Y(g4234),.A(g3793),.B(ttmp694));
OR2X1 OR_tmp696 (.Y(ttmp696),.A(g9569),.B(I15042));
OR2X1 OR_tmp697 (.Y(ttmp697),.A(g9512),.B(ttmp696));
NOR2X1 NOR_tmp698 (.Y(g9877),.A(g9536),.B(ttmp697));
NOR2X1 NOR2_87 (.Y(g5186),.A(g2047),.B(g4401));
NOR2X1 NOR2_88 (.Y(g9489),.A(g9052),.B(g9030));
OR2X1 OR_tmp699 (.Y(ttmp699),.A(g3485),.B(g2655));
OR2X1 OR_tmp700 (.Y(ttmp700),.A(g3077),.B(ttmp699));
NOR2X1 NOR_tmp701 (.Y(g4619),.A(g3491),.B(ttmp700));
NOR2X1 NOR2_89 (.Y(g10432),.A(g10350),.B(g3566));
NOR2X1 NOR2_90 (.Y(g5345),.A(g2754),.B(g4835));
NOR2X1 NOR2_91 (.Y(g5763),.A(g5350),.B(g5345));
NOR2X1 NOR2_92 (.Y(g10375),.A(g10288),.B(g3463));
OR2X1 OR_tmp702 (.Y(ttmp702),.A(g3784),.B(g2579));
OR2X1 OR_tmp703 (.Y(ttmp703),.A(g3292),.B(ttmp702));
NOR2X1 NOR_tmp704 (.Y(g4879),.A(g2593),.B(ttmp703));
NOR2X1 OR_tmp705 (.Y(ttmp705),.A(g3485),.B(g3479));
OR2X1 OR_tmp706 (.Y(ttmp706),.A(g3077),.B(ttmp705));
OR2X1 NOR_tmp707 (.Y(g4607),.A(g2669),.B(ttmp706));
NOR2X1 NOR2_93 (.Y(g10425),.A(g10293),.B(g4620));
OR2X1 NOR2_94 (.Y(g3107),.A(g2501),.B(g2499));
NOR2X1 NOR2_95 (.Y(g10322),.A(g9317),.B(g10272));
OR2X1 OR_tmp708 (.Y(ttmp708),.A(g3485),.B(g3479));
NOR2X1 OR_tmp709 (.Y(ttmp709),.A(g3077),.B(ttmp708));
NOR2X1 NOR_tmp710 (.Y(g4630),.A(g3491),.B(ttmp709));
NOR2X1 NOR2_96 (.Y(g10364),.A(g10327),.B(g3744));
NOR2X1 NOR2_97 (.Y(g9781),.A(g9392),.B(g9367));
endmodule
